// q_sys.v

// Generated using ACDS version 19.1 670

`timescale 1 ps / 1 ps
module q_sys (
		output wire        altpll_shift_c0_clk,                         //                     altpll_shift_c0.clk
		output wire        altpll_shift_locked_conduit_export,          //         altpll_shift_locked_conduit.export
		input  wire [8:0]  button_pio_external_connection_export,       //      button_pio_external_connection.export
		input  wire        clock_bridge_0_in_clk_clk,                   //               clock_bridge_0_in_clk.clk
		input  wire        ddr3_ram_pll_ref_clk_clk,                    //                ddr3_ram_pll_ref_clk.clk
		input  wire        debug_uart_external_connection_rxd,          //      debug_uart_external_connection.rxd
		output wire        debug_uart_external_connection_txd,          //                                    .txd
		output wire        enet_pll_c0_clk,                             //                         enet_pll_c0.clk
		output wire        enet_pll_c1_clk,                             //                         enet_pll_c1.clk
		output wire        enet_pll_c2_clk,                             //                         enet_pll_c2.clk
		output wire        enet_pll_c3_clk,                             //                         enet_pll_c3.clk
		output wire        enet_pll_c4_clk,                             //                         enet_pll_c4.clk
		output wire        enet_pll_locked_conduit_export,              //             enet_pll_locked_conduit.export
		output wire        eth_tse_mac_mdio_connection_mdc,             //         eth_tse_mac_mdio_connection.mdc
		input  wire        eth_tse_mac_mdio_connection_mdio_in,         //                                    .mdio_in
		output wire        eth_tse_mac_mdio_connection_mdio_out,        //                                    .mdio_out
		output wire        eth_tse_mac_mdio_connection_mdio_oen,        //                                    .mdio_oen
		input  wire [3:0]  eth_tse_mac_rgmii_connection_rgmii_in,       //        eth_tse_mac_rgmii_connection.rgmii_in
		output wire [3:0]  eth_tse_mac_rgmii_connection_rgmii_out,      //                                    .rgmii_out
		input  wire        eth_tse_mac_rgmii_connection_rx_control,     //                                    .rx_control
		output wire        eth_tse_mac_rgmii_connection_tx_control,     //                                    .tx_control
		input  wire        eth_tse_mac_status_connection_set_10,        //       eth_tse_mac_status_connection.set_10
		input  wire        eth_tse_mac_status_connection_set_1000,      //                                    .set_1000
		output wire        eth_tse_mac_status_connection_eth_mode,      //                                    .eth_mode
		output wire        eth_tse_mac_status_connection_ena_10,        //                                    .ena_10
		input  wire        eth_tse_pcs_mac_rx_clock_connection_clk,     // eth_tse_pcs_mac_rx_clock_connection.clk
		input  wire        eth_tse_pcs_mac_tx_clock_connection_clk,     // eth_tse_pcs_mac_tx_clock_connection.clk
		inout  wire [3:0]  ext_flash_flash_dataout_conduit_dataout,     //             ext_flash_flash_dataout.conduit_dataout
		output wire        ext_flash_flash_dclk_out_conduit_dclk_out,   //            ext_flash_flash_dclk_out.conduit_dclk_out
		output wire [0:0]  ext_flash_flash_ncs_conduit_ncs,             //                 ext_flash_flash_ncs.conduit_ncs
		output wire        frame_timer_export,                          //                         frame_timer.export
		output wire [7:0]  led_pio_external_connection_export,          //         led_pio_external_connection.export
		output wire        mem_if_ddr3_emif_0_status_local_init_done,   //           mem_if_ddr3_emif_0_status.local_init_done
		output wire        mem_if_ddr3_emif_0_status_local_cal_success, //                                    .local_cal_success
		output wire        mem_if_ddr3_emif_0_status_local_cal_fail,    //                                    .local_cal_fail
		input  wire        mem_resetn_in_reset_reset_n,                 //                 mem_resetn_in_reset.reset_n
		output wire [13:0] memory_mem_a,                                //                              memory.mem_a
		output wire [2:0]  memory_mem_ba,                               //                                    .mem_ba
		inout  wire [0:0]  memory_mem_ck,                               //                                    .mem_ck
		inout  wire [0:0]  memory_mem_ck_n,                             //                                    .mem_ck_n
		output wire [0:0]  memory_mem_cke,                              //                                    .mem_cke
		output wire [0:0]  memory_mem_cs_n,                             //                                    .mem_cs_n
		output wire [0:0]  memory_mem_dm,                               //                                    .mem_dm
		output wire [0:0]  memory_mem_ras_n,                            //                                    .mem_ras_n
		output wire [0:0]  memory_mem_cas_n,                            //                                    .mem_cas_n
		output wire [0:0]  memory_mem_we_n,                             //                                    .mem_we_n
		output wire        memory_mem_reset_n,                          //                                    .mem_reset_n
		inout  wire [7:0]  memory_mem_dq,                               //                                    .mem_dq
		inout  wire [0:0]  memory_mem_dqs,                              //                                    .mem_dqs
		inout  wire [0:0]  memory_mem_dqs_n,                            //                                    .mem_dqs_n
		output wire [0:0]  memory_mem_odt,                              //                                    .mem_odt
		input  wire        reset_reset_n,                               //                               reset.reset_n
		input  wire [4:0]  sensor_in_adc_data,                          //                              sensor.in_adc_data
		input  wire        sensor_in_trg,                               //                                    .in_trg
		output wire        sensor_out_adc_clk,                          //                                    .out_adc_clk
		output wire        sensor_out_adc_cnv,                          //                                    .out_adc_cnv
		output wire        sensor_out_sensor_clk,                       //                                    .out_sensor_clk
		output wire        sensor_out_sensor_gain,                      //                                    .out_sensor_gain
		output wire        sensor_out_sensor_rst,                       //                                    .out_sensor_rst
		output wire [7:0]  sensor_status_status_out,                    //                       sensor_status.status_out
		input  wire [7:0]  sensor_synchro_ext_input,                    //                      sensor_synchro.ext_input
		input  wire        sensor_synchro_serial_rx,                    //                                    .serial_rx
		output wire        sensor_synchro_serial_tx,                    //                                    .serial_tx
		input  wire        sys_clk_clk                                  //                             sys_clk.clk
	);

	wire         sensor_interface_data_out_valid;                        // sensor_interface:data_out_valid -> udp_generator:data_in_valid
	wire  [31:0] sensor_interface_data_out_data;                         // sensor_interface:data_out_data -> udp_generator:data_in_data
	wire         sensor_interface_data_out_ready;                        // udp_generator:data_in_ready -> sensor_interface:data_out_ready
	wire         sensor_interface_data_out_startofpacket;                // sensor_interface:data_out_startofpacket -> udp_generator:data_in_startofpacket
	wire         sensor_interface_data_out_endofpacket;                  // sensor_interface:data_out_endofpacket -> udp_generator:data_in_endofpacket
	wire   [1:0] sensor_interface_data_out_empty;                        // sensor_interface:data_out_empty -> udp_generator:data_in_empty
	wire         tx_multiplexer_out_valid;                               // tx_multiplexer:out_valid -> channel_adapter_0:in_valid
	wire  [31:0] tx_multiplexer_out_data;                                // tx_multiplexer:out_data -> channel_adapter_0:in_data
	wire         tx_multiplexer_out_ready;                               // channel_adapter_0:in_ready -> tx_multiplexer:out_ready
	wire         tx_multiplexer_out_channel;                             // tx_multiplexer:out_channel -> channel_adapter_0:in_channel
	wire         tx_multiplexer_out_startofpacket;                       // tx_multiplexer:out_startofpacket -> channel_adapter_0:in_startofpacket
	wire         tx_multiplexer_out_endofpacket;                         // tx_multiplexer:out_endofpacket -> channel_adapter_0:in_endofpacket
	wire         tx_multiplexer_out_error;                               // tx_multiplexer:out_error -> channel_adapter_0:in_error
	wire   [1:0] tx_multiplexer_out_empty;                               // tx_multiplexer:out_empty -> channel_adapter_0:in_empty
	wire         channel_adapter_0_out_valid;                            // channel_adapter_0:out_valid -> eth_tse:ff_tx_wren
	wire  [31:0] channel_adapter_0_out_data;                             // channel_adapter_0:out_data -> eth_tse:ff_tx_data
	wire         channel_adapter_0_out_ready;                            // eth_tse:ff_tx_rdy -> channel_adapter_0:out_ready
	wire         channel_adapter_0_out_startofpacket;                    // channel_adapter_0:out_startofpacket -> eth_tse:ff_tx_sop
	wire         channel_adapter_0_out_endofpacket;                      // channel_adapter_0:out_endofpacket -> eth_tse:ff_tx_eop
	wire         channel_adapter_0_out_error;                            // channel_adapter_0:out_error -> eth_tse:ff_tx_err
	wire   [1:0] channel_adapter_0_out_empty;                            // channel_adapter_0:out_empty -> eth_tse:ff_tx_mod
	wire         msgdma_tx_st_source_valid;                              // msgdma_tx:st_source_valid -> tx_multiplexer:in0_valid
	wire  [31:0] msgdma_tx_st_source_data;                               // msgdma_tx:st_source_data -> tx_multiplexer:in0_data
	wire         msgdma_tx_st_source_ready;                              // tx_multiplexer:in0_ready -> msgdma_tx:st_source_ready
	wire         msgdma_tx_st_source_startofpacket;                      // msgdma_tx:st_source_startofpacket -> tx_multiplexer:in0_startofpacket
	wire         msgdma_tx_st_source_endofpacket;                        // msgdma_tx:st_source_endofpacket -> tx_multiplexer:in0_endofpacket
	wire         msgdma_tx_st_source_error;                              // msgdma_tx:st_source_error -> tx_multiplexer:in0_error
	wire   [1:0] msgdma_tx_st_source_empty;                              // msgdma_tx:st_source_empty -> tx_multiplexer:in0_empty
	wire  [15:0] sensor_interface_calibration_ram_interface_readdata;    // mm_interconnect_0:sensor_interface_calibration_ram_interface_readdata -> sensor_interface:cali_fac
	wire         sensor_interface_calibration_ram_interface_waitrequest; // mm_interconnect_0:sensor_interface_calibration_ram_interface_waitrequest -> sensor_interface:waitrequest
	wire   [8:0] sensor_interface_calibration_ram_interface_address;     // sensor_interface:address -> mm_interconnect_0:sensor_interface_calibration_ram_interface_address
	wire         sensor_interface_calibration_ram_interface_read;        // sensor_interface:clken -> mm_interconnect_0:sensor_interface_calibration_ram_interface_read
	wire         mm_interconnect_0_calibration_ram_s2_chipselect;        // mm_interconnect_0:calibration_ram_s2_chipselect -> calibration_ram:chipselect2
	wire  [15:0] mm_interconnect_0_calibration_ram_s2_readdata;          // calibration_ram:readdata2 -> mm_interconnect_0:calibration_ram_s2_readdata
	wire   [8:0] mm_interconnect_0_calibration_ram_s2_address;           // mm_interconnect_0:calibration_ram_s2_address -> calibration_ram:address2
	wire   [1:0] mm_interconnect_0_calibration_ram_s2_byteenable;        // mm_interconnect_0:calibration_ram_s2_byteenable -> calibration_ram:byteenable2
	wire         mm_interconnect_0_calibration_ram_s2_write;             // mm_interconnect_0:calibration_ram_s2_write -> calibration_ram:write2
	wire  [15:0] mm_interconnect_0_calibration_ram_s2_writedata;         // mm_interconnect_0:calibration_ram_s2_writedata -> calibration_ram:writedata2
	wire         mm_interconnect_0_calibration_ram_s2_clken;             // mm_interconnect_0:calibration_ram_s2_clken -> calibration_ram:clken2
	wire  [31:0] cpu_data_master_readdata;                               // mm_interconnect_1:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                            // mm_interconnect_1:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                            // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_1:cpu_data_master_debugaccess
	wire  [28:0] cpu_data_master_address;                                // cpu:d_address -> mm_interconnect_1:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                             // cpu:d_byteenable -> mm_interconnect_1:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                   // cpu:d_read -> mm_interconnect_1:cpu_data_master_read
	wire         cpu_data_master_readdatavalid;                          // mm_interconnect_1:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	wire         cpu_data_master_write;                                  // cpu:d_write -> mm_interconnect_1:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                              // cpu:d_writedata -> mm_interconnect_1:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                        // mm_interconnect_1:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                     // mm_interconnect_1:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [28:0] cpu_instruction_master_address;                         // cpu:i_address -> mm_interconnect_1:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                            // cpu:i_read -> mm_interconnect_1:cpu_instruction_master_read
	wire         cpu_instruction_master_readdatavalid;                   // mm_interconnect_1:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire  [31:0] msgdma_tx_mm_read_readdata;                             // mm_interconnect_1:msgdma_tx_mm_read_readdata -> msgdma_tx:mm_read_readdata
	wire         msgdma_tx_mm_read_waitrequest;                          // mm_interconnect_1:msgdma_tx_mm_read_waitrequest -> msgdma_tx:mm_read_waitrequest
	wire  [27:0] msgdma_tx_mm_read_address;                              // msgdma_tx:mm_read_address -> mm_interconnect_1:msgdma_tx_mm_read_address
	wire         msgdma_tx_mm_read_read;                                 // msgdma_tx:mm_read_read -> mm_interconnect_1:msgdma_tx_mm_read_read
	wire   [3:0] msgdma_tx_mm_read_byteenable;                           // msgdma_tx:mm_read_byteenable -> mm_interconnect_1:msgdma_tx_mm_read_byteenable
	wire         msgdma_tx_mm_read_readdatavalid;                        // mm_interconnect_1:msgdma_tx_mm_read_readdatavalid -> msgdma_tx:mm_read_readdatavalid
	wire         msgdma_rx_mm_write_waitrequest;                         // mm_interconnect_1:msgdma_rx_mm_write_waitrequest -> msgdma_rx:mm_write_waitrequest
	wire  [27:0] msgdma_rx_mm_write_address;                             // msgdma_rx:mm_write_address -> mm_interconnect_1:msgdma_rx_mm_write_address
	wire   [3:0] msgdma_rx_mm_write_byteenable;                          // msgdma_rx:mm_write_byteenable -> mm_interconnect_1:msgdma_rx_mm_write_byteenable
	wire         msgdma_rx_mm_write_write;                               // msgdma_rx:mm_write_write -> mm_interconnect_1:msgdma_rx_mm_write_write
	wire  [31:0] msgdma_rx_mm_write_writedata;                           // msgdma_rx:mm_write_writedata -> mm_interconnect_1:msgdma_rx_mm_write_writedata
	wire  [31:0] msgdma_tx_descriptor_read_master_readdata;              // mm_interconnect_1:msgdma_tx_descriptor_read_master_readdata -> msgdma_tx:descriptor_read_master_readdata
	wire         msgdma_tx_descriptor_read_master_waitrequest;           // mm_interconnect_1:msgdma_tx_descriptor_read_master_waitrequest -> msgdma_tx:descriptor_read_master_waitrequest
	wire  [28:0] msgdma_tx_descriptor_read_master_address;               // msgdma_tx:descriptor_read_master_address -> mm_interconnect_1:msgdma_tx_descriptor_read_master_address
	wire         msgdma_tx_descriptor_read_master_read;                  // msgdma_tx:descriptor_read_master_read -> mm_interconnect_1:msgdma_tx_descriptor_read_master_read
	wire         msgdma_tx_descriptor_read_master_readdatavalid;         // mm_interconnect_1:msgdma_tx_descriptor_read_master_readdatavalid -> msgdma_tx:descriptor_read_master_readdatavalid
	wire  [31:0] msgdma_rx_descriptor_read_master_readdata;              // mm_interconnect_1:msgdma_rx_descriptor_read_master_readdata -> msgdma_rx:descriptor_read_master_readdata
	wire         msgdma_rx_descriptor_read_master_waitrequest;           // mm_interconnect_1:msgdma_rx_descriptor_read_master_waitrequest -> msgdma_rx:descriptor_read_master_waitrequest
	wire  [28:0] msgdma_rx_descriptor_read_master_address;               // msgdma_rx:descriptor_read_master_address -> mm_interconnect_1:msgdma_rx_descriptor_read_master_address
	wire         msgdma_rx_descriptor_read_master_read;                  // msgdma_rx:descriptor_read_master_read -> mm_interconnect_1:msgdma_rx_descriptor_read_master_read
	wire         msgdma_rx_descriptor_read_master_readdatavalid;         // mm_interconnect_1:msgdma_rx_descriptor_read_master_readdatavalid -> msgdma_rx:descriptor_read_master_readdatavalid
	wire         msgdma_tx_descriptor_write_master_waitrequest;          // mm_interconnect_1:msgdma_tx_descriptor_write_master_waitrequest -> msgdma_tx:descriptor_write_master_waitrequest
	wire  [28:0] msgdma_tx_descriptor_write_master_address;              // msgdma_tx:descriptor_write_master_address -> mm_interconnect_1:msgdma_tx_descriptor_write_master_address
	wire   [3:0] msgdma_tx_descriptor_write_master_byteenable;           // msgdma_tx:descriptor_write_master_byteenable -> mm_interconnect_1:msgdma_tx_descriptor_write_master_byteenable
	wire   [1:0] msgdma_tx_descriptor_write_master_response;             // mm_interconnect_1:msgdma_tx_descriptor_write_master_response -> msgdma_tx:descriptor_write_master_response
	wire         msgdma_tx_descriptor_write_master_write;                // msgdma_tx:descriptor_write_master_write -> mm_interconnect_1:msgdma_tx_descriptor_write_master_write
	wire  [31:0] msgdma_tx_descriptor_write_master_writedata;            // msgdma_tx:descriptor_write_master_writedata -> mm_interconnect_1:msgdma_tx_descriptor_write_master_writedata
	wire         msgdma_tx_descriptor_write_master_writeresponsevalid;   // mm_interconnect_1:msgdma_tx_descriptor_write_master_writeresponsevalid -> msgdma_tx:descriptor_write_master_writeresponsevalid
	wire         msgdma_rx_descriptor_write_master_waitrequest;          // mm_interconnect_1:msgdma_rx_descriptor_write_master_waitrequest -> msgdma_rx:descriptor_write_master_waitrequest
	wire  [28:0] msgdma_rx_descriptor_write_master_address;              // msgdma_rx:descriptor_write_master_address -> mm_interconnect_1:msgdma_rx_descriptor_write_master_address
	wire   [3:0] msgdma_rx_descriptor_write_master_byteenable;           // msgdma_rx:descriptor_write_master_byteenable -> mm_interconnect_1:msgdma_rx_descriptor_write_master_byteenable
	wire   [1:0] msgdma_rx_descriptor_write_master_response;             // mm_interconnect_1:msgdma_rx_descriptor_write_master_response -> msgdma_rx:descriptor_write_master_response
	wire         msgdma_rx_descriptor_write_master_write;                // msgdma_rx:descriptor_write_master_write -> mm_interconnect_1:msgdma_rx_descriptor_write_master_write
	wire  [31:0] msgdma_rx_descriptor_write_master_writedata;            // msgdma_rx:descriptor_write_master_writedata -> mm_interconnect_1:msgdma_rx_descriptor_write_master_writedata
	wire         msgdma_rx_descriptor_write_master_writeresponsevalid;   // mm_interconnect_1:msgdma_rx_descriptor_write_master_writeresponsevalid -> msgdma_rx:descriptor_write_master_writeresponsevalid
	wire         mm_interconnect_1_ddr3_ram_avl_beginbursttransfer;      // mm_interconnect_1:ddr3_ram_avl_beginbursttransfer -> ddr3_ram:avl_burstbegin
	wire  [31:0] mm_interconnect_1_ddr3_ram_avl_readdata;                // ddr3_ram:avl_rdata -> mm_interconnect_1:ddr3_ram_avl_readdata
	wire         mm_interconnect_1_ddr3_ram_avl_waitrequest;             // ddr3_ram:avl_ready -> mm_interconnect_1:ddr3_ram_avl_waitrequest
	wire  [24:0] mm_interconnect_1_ddr3_ram_avl_address;                 // mm_interconnect_1:ddr3_ram_avl_address -> ddr3_ram:avl_addr
	wire         mm_interconnect_1_ddr3_ram_avl_read;                    // mm_interconnect_1:ddr3_ram_avl_read -> ddr3_ram:avl_read_req
	wire   [3:0] mm_interconnect_1_ddr3_ram_avl_byteenable;              // mm_interconnect_1:ddr3_ram_avl_byteenable -> ddr3_ram:avl_be
	wire         mm_interconnect_1_ddr3_ram_avl_readdatavalid;           // ddr3_ram:avl_rdata_valid -> mm_interconnect_1:ddr3_ram_avl_readdatavalid
	wire         mm_interconnect_1_ddr3_ram_avl_write;                   // mm_interconnect_1:ddr3_ram_avl_write -> ddr3_ram:avl_write_req
	wire  [31:0] mm_interconnect_1_ddr3_ram_avl_writedata;               // mm_interconnect_1:ddr3_ram_avl_writedata -> ddr3_ram:avl_wdata
	wire   [2:0] mm_interconnect_1_ddr3_ram_avl_burstcount;              // mm_interconnect_1:ddr3_ram_avl_burstcount -> ddr3_ram:avl_size
	wire         ddr3_ram_afi_clk_clk;                                   // ddr3_ram:afi_clk -> [mm_interconnect_1:ddr3_ram_afi_clk_clk, rst_controller_006:clk]
	wire  [31:0] mm_interconnect_1_ext_flash_avl_csr_readdata;           // ext_flash:avl_csr_rddata -> mm_interconnect_1:ext_flash_avl_csr_readdata
	wire         mm_interconnect_1_ext_flash_avl_csr_waitrequest;        // ext_flash:avl_csr_waitrequest -> mm_interconnect_1:ext_flash_avl_csr_waitrequest
	wire   [2:0] mm_interconnect_1_ext_flash_avl_csr_address;            // mm_interconnect_1:ext_flash_avl_csr_address -> ext_flash:avl_csr_addr
	wire         mm_interconnect_1_ext_flash_avl_csr_read;               // mm_interconnect_1:ext_flash_avl_csr_read -> ext_flash:avl_csr_read
	wire         mm_interconnect_1_ext_flash_avl_csr_readdatavalid;      // ext_flash:avl_csr_rddata_valid -> mm_interconnect_1:ext_flash_avl_csr_readdatavalid
	wire         mm_interconnect_1_ext_flash_avl_csr_write;              // mm_interconnect_1:ext_flash_avl_csr_write -> ext_flash:avl_csr_write
	wire  [31:0] mm_interconnect_1_ext_flash_avl_csr_writedata;          // mm_interconnect_1:ext_flash_avl_csr_writedata -> ext_flash:avl_csr_wrdata
	wire  [31:0] mm_interconnect_1_ext_flash_avl_mem_readdata;           // ext_flash:avl_mem_rddata -> mm_interconnect_1:ext_flash_avl_mem_readdata
	wire         mm_interconnect_1_ext_flash_avl_mem_waitrequest;        // ext_flash:avl_mem_waitrequest -> mm_interconnect_1:ext_flash_avl_mem_waitrequest
	wire  [23:0] mm_interconnect_1_ext_flash_avl_mem_address;            // mm_interconnect_1:ext_flash_avl_mem_address -> ext_flash:avl_mem_addr
	wire         mm_interconnect_1_ext_flash_avl_mem_read;               // mm_interconnect_1:ext_flash_avl_mem_read -> ext_flash:avl_mem_read
	wire   [3:0] mm_interconnect_1_ext_flash_avl_mem_byteenable;         // mm_interconnect_1:ext_flash_avl_mem_byteenable -> ext_flash:avl_mem_byteenable
	wire         mm_interconnect_1_ext_flash_avl_mem_readdatavalid;      // ext_flash:avl_mem_rddata_valid -> mm_interconnect_1:ext_flash_avl_mem_readdatavalid
	wire         mm_interconnect_1_ext_flash_avl_mem_write;              // mm_interconnect_1:ext_flash_avl_mem_write -> ext_flash:avl_mem_write
	wire  [31:0] mm_interconnect_1_ext_flash_avl_mem_writedata;          // mm_interconnect_1:ext_flash_avl_mem_writedata -> ext_flash:avl_mem_wrdata
	wire   [6:0] mm_interconnect_1_ext_flash_avl_mem_burstcount;         // mm_interconnect_1:ext_flash_avl_mem_burstcount -> ext_flash:avl_mem_burstcount
	wire  [31:0] mm_interconnect_1_eth_tse_control_port_readdata;        // eth_tse:reg_data_out -> mm_interconnect_1:eth_tse_control_port_readdata
	wire         mm_interconnect_1_eth_tse_control_port_waitrequest;     // eth_tse:reg_busy -> mm_interconnect_1:eth_tse_control_port_waitrequest
	wire   [7:0] mm_interconnect_1_eth_tse_control_port_address;         // mm_interconnect_1:eth_tse_control_port_address -> eth_tse:reg_addr
	wire         mm_interconnect_1_eth_tse_control_port_read;            // mm_interconnect_1:eth_tse_control_port_read -> eth_tse:reg_rd
	wire         mm_interconnect_1_eth_tse_control_port_write;           // mm_interconnect_1:eth_tse_control_port_write -> eth_tse:reg_wr
	wire  [31:0] mm_interconnect_1_eth_tse_control_port_writedata;       // mm_interconnect_1:eth_tse_control_port_writedata -> eth_tse:reg_data_in
	wire  [31:0] mm_interconnect_1_sysid_control_slave_readdata;         // sysid:readdata -> mm_interconnect_1:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_1_sysid_control_slave_address;          // mm_interconnect_1:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_1_msgdma_tx_csr_readdata;               // msgdma_tx:csr_readdata -> mm_interconnect_1:msgdma_tx_csr_readdata
	wire   [2:0] mm_interconnect_1_msgdma_tx_csr_address;                // mm_interconnect_1:msgdma_tx_csr_address -> msgdma_tx:csr_address
	wire         mm_interconnect_1_msgdma_tx_csr_read;                   // mm_interconnect_1:msgdma_tx_csr_read -> msgdma_tx:csr_read
	wire   [3:0] mm_interconnect_1_msgdma_tx_csr_byteenable;             // mm_interconnect_1:msgdma_tx_csr_byteenable -> msgdma_tx:csr_byteenable
	wire         mm_interconnect_1_msgdma_tx_csr_write;                  // mm_interconnect_1:msgdma_tx_csr_write -> msgdma_tx:csr_write
	wire  [31:0] mm_interconnect_1_msgdma_tx_csr_writedata;              // mm_interconnect_1:msgdma_tx_csr_writedata -> msgdma_tx:csr_writedata
	wire  [31:0] mm_interconnect_1_msgdma_rx_csr_readdata;               // msgdma_rx:csr_readdata -> mm_interconnect_1:msgdma_rx_csr_readdata
	wire   [2:0] mm_interconnect_1_msgdma_rx_csr_address;                // mm_interconnect_1:msgdma_rx_csr_address -> msgdma_rx:csr_address
	wire         mm_interconnect_1_msgdma_rx_csr_read;                   // mm_interconnect_1:msgdma_rx_csr_read -> msgdma_rx:csr_read
	wire   [3:0] mm_interconnect_1_msgdma_rx_csr_byteenable;             // mm_interconnect_1:msgdma_rx_csr_byteenable -> msgdma_rx:csr_byteenable
	wire         mm_interconnect_1_msgdma_rx_csr_write;                  // mm_interconnect_1:msgdma_rx_csr_write -> msgdma_rx:csr_write
	wire  [31:0] mm_interconnect_1_msgdma_rx_csr_writedata;              // mm_interconnect_1:msgdma_rx_csr_writedata -> msgdma_rx:csr_writedata
	wire  [31:0] mm_interconnect_1_onchip_flash_csr_readdata;            // onchip_flash:avmm_csr_readdata -> mm_interconnect_1:onchip_flash_csr_readdata
	wire   [0:0] mm_interconnect_1_onchip_flash_csr_address;             // mm_interconnect_1:onchip_flash_csr_address -> onchip_flash:avmm_csr_addr
	wire         mm_interconnect_1_onchip_flash_csr_read;                // mm_interconnect_1:onchip_flash_csr_read -> onchip_flash:avmm_csr_read
	wire         mm_interconnect_1_onchip_flash_csr_write;               // mm_interconnect_1:onchip_flash_csr_write -> onchip_flash:avmm_csr_write
	wire  [31:0] mm_interconnect_1_onchip_flash_csr_writedata;           // mm_interconnect_1:onchip_flash_csr_writedata -> onchip_flash:avmm_csr_writedata
	wire  [31:0] mm_interconnect_1_udp_generator_csr_readdata;           // udp_generator:csr_readdata -> mm_interconnect_1:udp_generator_csr_readdata
	wire   [2:0] mm_interconnect_1_udp_generator_csr_address;            // mm_interconnect_1:udp_generator_csr_address -> udp_generator:csr_address
	wire         mm_interconnect_1_udp_generator_csr_read;               // mm_interconnect_1:udp_generator_csr_read -> udp_generator:csr_read
	wire   [3:0] mm_interconnect_1_udp_generator_csr_byteenable;         // mm_interconnect_1:udp_generator_csr_byteenable -> udp_generator:csr_byteenable
	wire         mm_interconnect_1_udp_generator_csr_write;              // mm_interconnect_1:udp_generator_csr_write -> udp_generator:csr_write
	wire  [31:0] mm_interconnect_1_udp_generator_csr_writedata;          // mm_interconnect_1:udp_generator_csr_writedata -> udp_generator:csr_writedata
	wire  [31:0] mm_interconnect_1_sensor_interface_csr_readdata;        // sensor_interface:csr_readdata -> mm_interconnect_1:sensor_interface_csr_readdata
	wire   [1:0] mm_interconnect_1_sensor_interface_csr_address;         // mm_interconnect_1:sensor_interface_csr_address -> sensor_interface:csr_address
	wire         mm_interconnect_1_sensor_interface_csr_read;            // mm_interconnect_1:sensor_interface_csr_read -> sensor_interface:csr_read
	wire   [3:0] mm_interconnect_1_sensor_interface_csr_byteenable;      // mm_interconnect_1:sensor_interface_csr_byteenable -> sensor_interface:csr_byteenable
	wire         mm_interconnect_1_sensor_interface_csr_write;           // mm_interconnect_1:sensor_interface_csr_write -> sensor_interface:csr_write
	wire  [31:0] mm_interconnect_1_sensor_interface_csr_writedata;       // mm_interconnect_1:sensor_interface_csr_writedata -> sensor_interface:csr_writedata
	wire  [31:0] mm_interconnect_1_onchip_flash_data_readdata;           // onchip_flash:avmm_data_readdata -> mm_interconnect_1:onchip_flash_data_readdata
	wire         mm_interconnect_1_onchip_flash_data_waitrequest;        // onchip_flash:avmm_data_waitrequest -> mm_interconnect_1:onchip_flash_data_waitrequest
	wire  [18:0] mm_interconnect_1_onchip_flash_data_address;            // mm_interconnect_1:onchip_flash_data_address -> onchip_flash:avmm_data_addr
	wire         mm_interconnect_1_onchip_flash_data_read;               // mm_interconnect_1:onchip_flash_data_read -> onchip_flash:avmm_data_read
	wire         mm_interconnect_1_onchip_flash_data_readdatavalid;      // onchip_flash:avmm_data_readdatavalid -> mm_interconnect_1:onchip_flash_data_readdatavalid
	wire         mm_interconnect_1_onchip_flash_data_write;              // mm_interconnect_1:onchip_flash_data_write -> onchip_flash:avmm_data_write
	wire  [31:0] mm_interconnect_1_onchip_flash_data_writedata;          // mm_interconnect_1:onchip_flash_data_writedata -> onchip_flash:avmm_data_writedata
	wire   [3:0] mm_interconnect_1_onchip_flash_data_burstcount;         // mm_interconnect_1:onchip_flash_data_burstcount -> onchip_flash:avmm_data_burstcount
	wire  [31:0] mm_interconnect_1_cpu_debug_mem_slave_readdata;         // cpu:debug_mem_slave_readdata -> mm_interconnect_1:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_1_cpu_debug_mem_slave_waitrequest;      // cpu:debug_mem_slave_waitrequest -> mm_interconnect_1:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_1_cpu_debug_mem_slave_debugaccess;      // mm_interconnect_1:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_1_cpu_debug_mem_slave_address;          // mm_interconnect_1:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_1_cpu_debug_mem_slave_read;             // mm_interconnect_1:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_1_cpu_debug_mem_slave_byteenable;       // mm_interconnect_1:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_1_cpu_debug_mem_slave_write;            // mm_interconnect_1:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_1_cpu_debug_mem_slave_writedata;        // mm_interconnect_1:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_1_msgdma_tx_prefetcher_csr_readdata;    // msgdma_tx:prefetcher_csr_readdata -> mm_interconnect_1:msgdma_tx_prefetcher_csr_readdata
	wire   [2:0] mm_interconnect_1_msgdma_tx_prefetcher_csr_address;     // mm_interconnect_1:msgdma_tx_prefetcher_csr_address -> msgdma_tx:prefetcher_csr_address
	wire         mm_interconnect_1_msgdma_tx_prefetcher_csr_read;        // mm_interconnect_1:msgdma_tx_prefetcher_csr_read -> msgdma_tx:prefetcher_csr_read
	wire         mm_interconnect_1_msgdma_tx_prefetcher_csr_write;       // mm_interconnect_1:msgdma_tx_prefetcher_csr_write -> msgdma_tx:prefetcher_csr_write
	wire  [31:0] mm_interconnect_1_msgdma_tx_prefetcher_csr_writedata;   // mm_interconnect_1:msgdma_tx_prefetcher_csr_writedata -> msgdma_tx:prefetcher_csr_writedata
	wire  [31:0] mm_interconnect_1_msgdma_rx_prefetcher_csr_readdata;    // msgdma_rx:prefetcher_csr_readdata -> mm_interconnect_1:msgdma_rx_prefetcher_csr_readdata
	wire   [2:0] mm_interconnect_1_msgdma_rx_prefetcher_csr_address;     // mm_interconnect_1:msgdma_rx_prefetcher_csr_address -> msgdma_rx:prefetcher_csr_address
	wire         mm_interconnect_1_msgdma_rx_prefetcher_csr_read;        // mm_interconnect_1:msgdma_rx_prefetcher_csr_read -> msgdma_rx:prefetcher_csr_read
	wire         mm_interconnect_1_msgdma_rx_prefetcher_csr_write;       // mm_interconnect_1:msgdma_rx_prefetcher_csr_write -> msgdma_rx:prefetcher_csr_write
	wire  [31:0] mm_interconnect_1_msgdma_rx_prefetcher_csr_writedata;   // mm_interconnect_1:msgdma_rx_prefetcher_csr_writedata -> msgdma_rx:prefetcher_csr_writedata
	wire         mm_interconnect_1_descriptor_memory_s1_chipselect;      // mm_interconnect_1:descriptor_memory_s1_chipselect -> descriptor_memory:chipselect
	wire  [31:0] mm_interconnect_1_descriptor_memory_s1_readdata;        // descriptor_memory:readdata -> mm_interconnect_1:descriptor_memory_s1_readdata
	wire  [10:0] mm_interconnect_1_descriptor_memory_s1_address;         // mm_interconnect_1:descriptor_memory_s1_address -> descriptor_memory:address
	wire   [3:0] mm_interconnect_1_descriptor_memory_s1_byteenable;      // mm_interconnect_1:descriptor_memory_s1_byteenable -> descriptor_memory:byteenable
	wire         mm_interconnect_1_descriptor_memory_s1_write;           // mm_interconnect_1:descriptor_memory_s1_write -> descriptor_memory:write
	wire  [31:0] mm_interconnect_1_descriptor_memory_s1_writedata;       // mm_interconnect_1:descriptor_memory_s1_writedata -> descriptor_memory:writedata
	wire         mm_interconnect_1_descriptor_memory_s1_clken;           // mm_interconnect_1:descriptor_memory_s1_clken -> descriptor_memory:clken
	wire         mm_interconnect_1_sys_clk_timer_s1_chipselect;          // mm_interconnect_1:sys_clk_timer_s1_chipselect -> sys_clk_timer:chipselect
	wire  [15:0] mm_interconnect_1_sys_clk_timer_s1_readdata;            // sys_clk_timer:readdata -> mm_interconnect_1:sys_clk_timer_s1_readdata
	wire   [2:0] mm_interconnect_1_sys_clk_timer_s1_address;             // mm_interconnect_1:sys_clk_timer_s1_address -> sys_clk_timer:address
	wire         mm_interconnect_1_sys_clk_timer_s1_write;               // mm_interconnect_1:sys_clk_timer_s1_write -> sys_clk_timer:write_n
	wire  [15:0] mm_interconnect_1_sys_clk_timer_s1_writedata;           // mm_interconnect_1:sys_clk_timer_s1_writedata -> sys_clk_timer:writedata
	wire         mm_interconnect_1_output_pio_s1_chipselect;             // mm_interconnect_1:output_pio_s1_chipselect -> output_pio:chipselect
	wire  [31:0] mm_interconnect_1_output_pio_s1_readdata;               // output_pio:readdata -> mm_interconnect_1:output_pio_s1_readdata
	wire   [2:0] mm_interconnect_1_output_pio_s1_address;                // mm_interconnect_1:output_pio_s1_address -> output_pio:address
	wire         mm_interconnect_1_output_pio_s1_write;                  // mm_interconnect_1:output_pio_s1_write -> output_pio:write_n
	wire  [31:0] mm_interconnect_1_output_pio_s1_writedata;              // mm_interconnect_1:output_pio_s1_writedata -> output_pio:writedata
	wire  [31:0] mm_interconnect_1_button_pio_s1_readdata;               // button_pio:readdata -> mm_interconnect_1:button_pio_s1_readdata
	wire   [1:0] mm_interconnect_1_button_pio_s1_address;                // mm_interconnect_1:button_pio_s1_address -> button_pio:address
	wire         mm_interconnect_1_debug_uart_s1_chipselect;             // mm_interconnect_1:debug_uart_s1_chipselect -> debug_uart:chipselect
	wire  [15:0] mm_interconnect_1_debug_uart_s1_readdata;               // debug_uart:readdata -> mm_interconnect_1:debug_uart_s1_readdata
	wire   [2:0] mm_interconnect_1_debug_uart_s1_address;                // mm_interconnect_1:debug_uart_s1_address -> debug_uart:address
	wire         mm_interconnect_1_debug_uart_s1_read;                   // mm_interconnect_1:debug_uart_s1_read -> debug_uart:read_n
	wire         mm_interconnect_1_debug_uart_s1_begintransfer;          // mm_interconnect_1:debug_uart_s1_begintransfer -> debug_uart:begintransfer
	wire         mm_interconnect_1_debug_uart_s1_write;                  // mm_interconnect_1:debug_uart_s1_write -> debug_uart:write_n
	wire  [15:0] mm_interconnect_1_debug_uart_s1_writedata;              // mm_interconnect_1:debug_uart_s1_writedata -> debug_uart:writedata
	wire         mm_interconnect_1_frame_timer_s1_chipselect;            // mm_interconnect_1:frame_timer_s1_chipselect -> frame_timer:chipselect
	wire  [15:0] mm_interconnect_1_frame_timer_s1_readdata;              // frame_timer:readdata -> mm_interconnect_1:frame_timer_s1_readdata
	wire   [2:0] mm_interconnect_1_frame_timer_s1_address;               // mm_interconnect_1:frame_timer_s1_address -> frame_timer:address
	wire         mm_interconnect_1_frame_timer_s1_write;                 // mm_interconnect_1:frame_timer_s1_write -> frame_timer:write_n
	wire  [15:0] mm_interconnect_1_frame_timer_s1_writedata;             // mm_interconnect_1:frame_timer_s1_writedata -> frame_timer:writedata
	wire         mm_interconnect_1_calibration_ram_s1_chipselect;        // mm_interconnect_1:calibration_ram_s1_chipselect -> calibration_ram:chipselect
	wire  [15:0] mm_interconnect_1_calibration_ram_s1_readdata;          // calibration_ram:readdata -> mm_interconnect_1:calibration_ram_s1_readdata
	wire   [8:0] mm_interconnect_1_calibration_ram_s1_address;           // mm_interconnect_1:calibration_ram_s1_address -> calibration_ram:address
	wire   [1:0] mm_interconnect_1_calibration_ram_s1_byteenable;        // mm_interconnect_1:calibration_ram_s1_byteenable -> calibration_ram:byteenable
	wire         mm_interconnect_1_calibration_ram_s1_write;             // mm_interconnect_1:calibration_ram_s1_write -> calibration_ram:write
	wire  [15:0] mm_interconnect_1_calibration_ram_s1_writedata;         // mm_interconnect_1:calibration_ram_s1_writedata -> calibration_ram:writedata
	wire         mm_interconnect_1_calibration_ram_s1_clken;             // mm_interconnect_1:calibration_ram_s1_clken -> calibration_ram:clken
	wire         irq_mapper_receiver0_irq;                               // msgdma_tx:csr_irq_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                               // msgdma_rx:csr_irq_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver3_irq;                               // sys_clk_timer:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                               // debug_uart:irq -> irq_mapper:receiver4_irq
	wire  [31:0] cpu_irq_irq;                                            // irq_mapper:sender_irq -> cpu:irq
	wire         irq_mapper_receiver2_irq;                               // irq_synchronizer:sender_irq -> irq_mapper:receiver2_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                          // ext_flash:irq -> irq_synchronizer:receiver_irq
	wire         udp_generator_data_out_valid;                           // udp_generator:data_out_valid -> avalon_st_adapter:in_0_valid
	wire  [31:0] udp_generator_data_out_data;                            // udp_generator:data_out_data -> avalon_st_adapter:in_0_data
	wire         udp_generator_data_out_ready;                           // avalon_st_adapter:in_0_ready -> udp_generator:data_out_ready
	wire         udp_generator_data_out_startofpacket;                   // udp_generator:data_out_startofpacket -> avalon_st_adapter:in_0_startofpacket
	wire         udp_generator_data_out_endofpacket;                     // udp_generator:data_out_endofpacket -> avalon_st_adapter:in_0_endofpacket
	wire   [1:0] udp_generator_data_out_empty;                           // udp_generator:data_out_empty -> avalon_st_adapter:in_0_empty
	wire         avalon_st_adapter_out_0_valid;                          // avalon_st_adapter:out_0_valid -> tx_multiplexer:in1_valid
	wire  [31:0] avalon_st_adapter_out_0_data;                           // avalon_st_adapter:out_0_data -> tx_multiplexer:in1_data
	wire         avalon_st_adapter_out_0_ready;                          // tx_multiplexer:in1_ready -> avalon_st_adapter:out_0_ready
	wire         avalon_st_adapter_out_0_startofpacket;                  // avalon_st_adapter:out_0_startofpacket -> tx_multiplexer:in1_startofpacket
	wire         avalon_st_adapter_out_0_endofpacket;                    // avalon_st_adapter:out_0_endofpacket -> tx_multiplexer:in1_endofpacket
	wire   [0:0] avalon_st_adapter_out_0_error;                          // avalon_st_adapter:out_0_error -> tx_multiplexer:in1_error
	wire   [1:0] avalon_st_adapter_out_0_empty;                          // avalon_st_adapter:out_0_empty -> tx_multiplexer:in1_empty
	wire         eth_tse_receive_valid;                                  // eth_tse:ff_rx_dval -> avalon_st_adapter_001:in_0_valid
	wire  [31:0] eth_tse_receive_data;                                   // eth_tse:ff_rx_data -> avalon_st_adapter_001:in_0_data
	wire         eth_tse_receive_ready;                                  // avalon_st_adapter_001:in_0_ready -> eth_tse:ff_rx_rdy
	wire         eth_tse_receive_startofpacket;                          // eth_tse:ff_rx_sop -> avalon_st_adapter_001:in_0_startofpacket
	wire         eth_tse_receive_endofpacket;                            // eth_tse:ff_rx_eop -> avalon_st_adapter_001:in_0_endofpacket
	wire   [5:0] eth_tse_receive_error;                                  // eth_tse:rx_err -> avalon_st_adapter_001:in_0_error
	wire   [1:0] eth_tse_receive_empty;                                  // eth_tse:ff_rx_mod -> avalon_st_adapter_001:in_0_empty
	wire         avalon_st_adapter_001_out_0_valid;                      // avalon_st_adapter_001:out_0_valid -> msgdma_rx:st_sink_valid
	wire  [31:0] avalon_st_adapter_001_out_0_data;                       // avalon_st_adapter_001:out_0_data -> msgdma_rx:st_sink_data
	wire         avalon_st_adapter_001_out_0_ready;                      // msgdma_rx:st_sink_ready -> avalon_st_adapter_001:out_0_ready
	wire         avalon_st_adapter_001_out_0_startofpacket;              // avalon_st_adapter_001:out_0_startofpacket -> msgdma_rx:st_sink_startofpacket
	wire         avalon_st_adapter_001_out_0_endofpacket;                // avalon_st_adapter_001:out_0_endofpacket -> msgdma_rx:st_sink_endofpacket
	wire   [5:0] avalon_st_adapter_001_out_0_error;                      // avalon_st_adapter_001:out_0_error -> msgdma_rx:st_sink_error
	wire   [1:0] avalon_st_adapter_001_out_0_empty;                      // avalon_st_adapter_001:out_0_empty -> msgdma_rx:st_sink_empty
	wire         rst_controller_reset_out_reset;                         // rst_controller:reset_out -> [altpll_shift:reset, enet_pll:reset]
	wire         rst_controller_001_reset_out_reset;                     // rst_controller_001:reset_out -> [avalon_st_adapter:in_rst_0_reset, button_pio:reset_n, calibration_ram:reset, calibration_ram:reset2, channel_adapter_0:reset_n, cpu:reset_n, debug_uart:reset_n, frame_timer:reset_n, irq_mapper:reset, irq_synchronizer:sender_reset, mm_interconnect_0:sensor_interface_rst_reset_bridge_in_reset_reset, mm_interconnect_1:cpu_reset_reset_bridge_in_reset_reset, msgdma_rx:reset_n_reset_n, msgdma_tx:reset_n_reset_n, onchip_flash:reset_n, rst_translator:in_reset, sensor_interface:rst_reset, tx_multiplexer:reset_n, udp_generator:rst_reset]
	wire         rst_controller_001_reset_out_reset_req;                 // rst_controller_001:reset_req -> [cpu:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_002_reset_out_reset;                     // rst_controller_002:reset_out -> ddr3_ram:global_reset_n
	wire         cpu_debug_reset_request_reset;                          // cpu:debug_reset_request -> [rst_controller_002:reset_in0, rst_controller_003:reset_in0, rst_controller_004:reset_in1, rst_controller_005:reset_in1, rst_controller_006:reset_in0]
	wire         rst_controller_003_reset_out_reset;                     // rst_controller_003:reset_out -> ddr3_ram:soft_reset_n
	wire         rst_controller_004_reset_out_reset;                     // rst_controller_004:reset_out -> [avalon_st_adapter_001:in_rst_0_reset, descriptor_memory:reset, eth_tse:reset, mm_interconnect_1:eth_tse_reset_connection_reset_bridge_in_reset_reset, output_pio:reset_n, rst_translator_001:in_reset, sys_clk_timer:reset_n, sysid:reset_n]
	wire         rst_controller_004_reset_out_reset_req;                 // rst_controller_004:reset_req -> [descriptor_memory:reset_req, rst_translator_001:reset_req_in]
	wire         rst_controller_005_reset_out_reset;                     // rst_controller_005:reset_out -> [ext_flash:reset_n, irq_synchronizer:receiver_reset, mm_interconnect_1:ext_flash_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_006_reset_out_reset;                     // rst_controller_006:reset_out -> [mm_interconnect_1:ddr3_ram_avl_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_1:ddr3_ram_soft_reset_reset_bridge_in_reset_reset]

	q_sys_altpll_shift altpll_shift (
		.clk                (sys_clk_clk),                        //       inclk_interface.clk
		.reset              (rst_controller_reset_out_reset),     // inclk_interface_reset.reset
		.read               (),                                   //             pll_slave.read
		.write              (),                                   //                      .write
		.address            (),                                   //                      .address
		.readdata           (),                                   //                      .readdata
		.writedata          (),                                   //                      .writedata
		.c0                 (altpll_shift_c0_clk),                //                    c0.clk
		.areset             (),                                   //        areset_conduit.export
		.locked             (altpll_shift_locked_conduit_export), //        locked_conduit.export
		.scandone           (),                                   //           (terminated)
		.scandataout        (),                                   //           (terminated)
		.c3                 (),                                   //           (terminated)
		.c4                 (),                                   //           (terminated)
		.phasecounterselect (3'b000),                             //           (terminated)
		.phaseupdown        (1'b0),                               //           (terminated)
		.phasestep          (1'b0),                               //           (terminated)
		.scanclk            (1'b0),                               //           (terminated)
		.scanclkena         (1'b0),                               //           (terminated)
		.scandata           (1'b0),                               //           (terminated)
		.configupdate       (1'b0),                               //           (terminated)
		.c1                 (),                                   //           (terminated)
		.c2                 (),                                   //           (terminated)
		.phasedone          ()                                    //           (terminated)
	);

	q_sys_button_pio button_pio (
		.clk      (sys_clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_1_button_pio_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_button_pio_s1_readdata), //                    .readdata
		.in_port  (button_pio_external_connection_export)     // external_connection.export
	);

	q_sys_calibration_ram calibration_ram (
		.clk         (sys_clk_clk),                                     //   clk1.clk
		.address     (mm_interconnect_1_calibration_ram_s1_address),    //     s1.address
		.clken       (mm_interconnect_1_calibration_ram_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_1_calibration_ram_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_1_calibration_ram_s1_write),      //       .write
		.readdata    (mm_interconnect_1_calibration_ram_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_1_calibration_ram_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_1_calibration_ram_s1_byteenable), //       .byteenable
		.reset       (rst_controller_001_reset_out_reset),              // reset1.reset
		.address2    (mm_interconnect_0_calibration_ram_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_calibration_ram_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_calibration_ram_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_calibration_ram_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_calibration_ram_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_calibration_ram_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_calibration_ram_s2_byteenable), //       .byteenable
		.clk2        (sys_clk_clk),                                     //   clk2.clk
		.reset2      (rst_controller_001_reset_out_reset),              // reset2.reset
		.reset_req   (1'b0),                                            // (terminated)
		.freeze      (1'b0),                                            // (terminated)
		.reset_req2  (1'b0)                                             // (terminated)
	);

	q_sys_channel_adapter_0 channel_adapter_0 (
		.clk               (sys_clk_clk),                         //   clk.clk
		.reset_n           (~rst_controller_001_reset_out_reset), // reset.reset_n
		.in_data           (tx_multiplexer_out_data),             //    in.data
		.in_valid          (tx_multiplexer_out_valid),            //      .valid
		.in_ready          (tx_multiplexer_out_ready),            //      .ready
		.in_startofpacket  (tx_multiplexer_out_startofpacket),    //      .startofpacket
		.in_endofpacket    (tx_multiplexer_out_endofpacket),      //      .endofpacket
		.in_empty          (tx_multiplexer_out_empty),            //      .empty
		.in_error          (tx_multiplexer_out_error),            //      .error
		.in_channel        (tx_multiplexer_out_channel),          //      .channel
		.out_data          (channel_adapter_0_out_data),          //   out.data
		.out_valid         (channel_adapter_0_out_valid),         //      .valid
		.out_ready         (channel_adapter_0_out_ready),         //      .ready
		.out_startofpacket (channel_adapter_0_out_startofpacket), //      .startofpacket
		.out_endofpacket   (channel_adapter_0_out_endofpacket),   //      .endofpacket
		.out_empty         (channel_adapter_0_out_empty),         //      .empty
		.out_error         (channel_adapter_0_out_error)          //      .error
	);

	q_sys_cpu cpu (
		.clk                                 (sys_clk_clk),                                       //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),               //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),            //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (cpu_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_1_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_1_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_1_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_1_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_1_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_1_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_1_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_1_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	q_sys_ddr3_ram ddr3_ram (
		.pll_ref_clk        (ddr3_ram_pll_ref_clk_clk),                          //      pll_ref_clk.clk
		.global_reset_n     (~rst_controller_002_reset_out_reset),               //     global_reset.reset_n
		.soft_reset_n       (~rst_controller_003_reset_out_reset),               //       soft_reset.reset_n
		.afi_clk            (ddr3_ram_afi_clk_clk),                              //          afi_clk.clk
		.afi_half_clk       (),                                                  //     afi_half_clk.clk
		.afi_reset_n        (),                                                  //        afi_reset.reset_n
		.afi_reset_export_n (),                                                  // afi_reset_export.reset_n
		.mem_a              (memory_mem_a),                                      //           memory.mem_a
		.mem_ba             (memory_mem_ba),                                     //                 .mem_ba
		.mem_ck             (memory_mem_ck),                                     //                 .mem_ck
		.mem_ck_n           (memory_mem_ck_n),                                   //                 .mem_ck_n
		.mem_cke            (memory_mem_cke),                                    //                 .mem_cke
		.mem_cs_n           (memory_mem_cs_n),                                   //                 .mem_cs_n
		.mem_dm             (memory_mem_dm),                                     //                 .mem_dm
		.mem_ras_n          (memory_mem_ras_n),                                  //                 .mem_ras_n
		.mem_cas_n          (memory_mem_cas_n),                                  //                 .mem_cas_n
		.mem_we_n           (memory_mem_we_n),                                   //                 .mem_we_n
		.mem_reset_n        (memory_mem_reset_n),                                //                 .mem_reset_n
		.mem_dq             (memory_mem_dq),                                     //                 .mem_dq
		.mem_dqs            (memory_mem_dqs),                                    //                 .mem_dqs
		.mem_dqs_n          (memory_mem_dqs_n),                                  //                 .mem_dqs_n
		.mem_odt            (memory_mem_odt),                                    //                 .mem_odt
		.avl_ready          (mm_interconnect_1_ddr3_ram_avl_waitrequest),        //              avl.waitrequest_n
		.avl_burstbegin     (mm_interconnect_1_ddr3_ram_avl_beginbursttransfer), //                 .beginbursttransfer
		.avl_addr           (mm_interconnect_1_ddr3_ram_avl_address),            //                 .address
		.avl_rdata_valid    (mm_interconnect_1_ddr3_ram_avl_readdatavalid),      //                 .readdatavalid
		.avl_rdata          (mm_interconnect_1_ddr3_ram_avl_readdata),           //                 .readdata
		.avl_wdata          (mm_interconnect_1_ddr3_ram_avl_writedata),          //                 .writedata
		.avl_be             (mm_interconnect_1_ddr3_ram_avl_byteenable),         //                 .byteenable
		.avl_read_req       (mm_interconnect_1_ddr3_ram_avl_read),               //                 .read
		.avl_write_req      (mm_interconnect_1_ddr3_ram_avl_write),              //                 .write
		.avl_size           (mm_interconnect_1_ddr3_ram_avl_burstcount),         //                 .burstcount
		.local_init_done    (mem_if_ddr3_emif_0_status_local_init_done),         //           status.local_init_done
		.local_cal_success  (mem_if_ddr3_emif_0_status_local_cal_success),       //                 .local_cal_success
		.local_cal_fail     (mem_if_ddr3_emif_0_status_local_cal_fail),          //                 .local_cal_fail
		.pll_mem_clk        (),                                                  //      pll_sharing.pll_mem_clk
		.pll_write_clk      (),                                                  //                 .pll_write_clk
		.pll_locked         (),                                                  //                 .pll_locked
		.pll_capture0_clk   (),                                                  //                 .pll_capture0_clk
		.pll_capture1_clk   ()                                                   //                 .pll_capture1_clk
	);

	q_sys_debug_uart debug_uart (
		.clk           (sys_clk_clk),                                   //                 clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),           //               reset.reset_n
		.address       (mm_interconnect_1_debug_uart_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_1_debug_uart_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_1_debug_uart_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_1_debug_uart_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_1_debug_uart_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_1_debug_uart_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_1_debug_uart_s1_readdata),      //                    .readdata
		.rxd           (debug_uart_external_connection_rxd),            // external_connection.export
		.txd           (debug_uart_external_connection_txd),            //                    .export
		.irq           (irq_mapper_receiver4_irq)                       //                 irq.irq
	);

	q_sys_descriptor_memory descriptor_memory (
		.clk        (sys_clk_clk),                                       //   clk1.clk
		.address    (mm_interconnect_1_descriptor_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_1_descriptor_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_1_descriptor_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_1_descriptor_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_1_descriptor_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_1_descriptor_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_1_descriptor_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_004_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_004_reset_out_reset_req),            //       .reset_req
		.freeze     (1'b0)                                               // (terminated)
	);

	q_sys_enet_pll enet_pll (
		.clk                (sys_clk_clk),                    //       inclk_interface.clk
		.reset              (rst_controller_reset_out_reset), // inclk_interface_reset.reset
		.read               (),                               //             pll_slave.read
		.write              (),                               //                      .write
		.address            (),                               //                      .address
		.readdata           (),                               //                      .readdata
		.writedata          (),                               //                      .writedata
		.c0                 (enet_pll_c0_clk),                //                    c0.clk
		.c1                 (enet_pll_c1_clk),                //                    c1.clk
		.c2                 (enet_pll_c2_clk),                //                    c2.clk
		.c3                 (enet_pll_c3_clk),                //                    c3.clk
		.c4                 (enet_pll_c4_clk),                //                    c4.clk
		.locked             (enet_pll_locked_conduit_export), //        locked_conduit.export
		.scandone           (),                               //           (terminated)
		.scandataout        (),                               //           (terminated)
		.phasecounterselect (3'b000),                         //           (terminated)
		.phaseupdown        (1'b0),                           //           (terminated)
		.phasestep          (1'b0),                           //           (terminated)
		.scanclk            (1'b0),                           //           (terminated)
		.scanclkena         (1'b0),                           //           (terminated)
		.scandata           (1'b0),                           //           (terminated)
		.configupdate       (1'b0),                           //           (terminated)
		.areset             (1'b0),                           //           (terminated)
		.phasedone          ()                                //           (terminated)
	);

	q_sys_eth_tse eth_tse (
		.clk           (sys_clk_clk),                                        // control_port_clock_connection.clk
		.reset         (rst_controller_004_reset_out_reset),                 //              reset_connection.reset
		.reg_addr      (mm_interconnect_1_eth_tse_control_port_address),     //                  control_port.address
		.reg_data_out  (mm_interconnect_1_eth_tse_control_port_readdata),    //                              .readdata
		.reg_rd        (mm_interconnect_1_eth_tse_control_port_read),        //                              .read
		.reg_data_in   (mm_interconnect_1_eth_tse_control_port_writedata),   //                              .writedata
		.reg_wr        (mm_interconnect_1_eth_tse_control_port_write),       //                              .write
		.reg_busy      (mm_interconnect_1_eth_tse_control_port_waitrequest), //                              .waitrequest
		.tx_clk        (eth_tse_pcs_mac_tx_clock_connection_clk),            //   pcs_mac_tx_clock_connection.clk
		.rx_clk        (eth_tse_pcs_mac_rx_clock_connection_clk),            //   pcs_mac_rx_clock_connection.clk
		.set_10        (eth_tse_mac_status_connection_set_10),               //         mac_status_connection.set_10
		.set_1000      (eth_tse_mac_status_connection_set_1000),             //                              .set_1000
		.eth_mode      (eth_tse_mac_status_connection_eth_mode),             //                              .eth_mode
		.ena_10        (eth_tse_mac_status_connection_ena_10),               //                              .ena_10
		.rgmii_in      (eth_tse_mac_rgmii_connection_rgmii_in),              //          mac_rgmii_connection.rgmii_in
		.rgmii_out     (eth_tse_mac_rgmii_connection_rgmii_out),             //                              .rgmii_out
		.rx_control    (eth_tse_mac_rgmii_connection_rx_control),            //                              .rx_control
		.tx_control    (eth_tse_mac_rgmii_connection_tx_control),            //                              .tx_control
		.ff_rx_clk     (sys_clk_clk),                                        //      receive_clock_connection.clk
		.ff_tx_clk     (sys_clk_clk),                                        //     transmit_clock_connection.clk
		.ff_rx_data    (eth_tse_receive_data),                               //                       receive.data
		.ff_rx_eop     (eth_tse_receive_endofpacket),                        //                              .endofpacket
		.rx_err        (eth_tse_receive_error),                              //                              .error
		.ff_rx_mod     (eth_tse_receive_empty),                              //                              .empty
		.ff_rx_rdy     (eth_tse_receive_ready),                              //                              .ready
		.ff_rx_sop     (eth_tse_receive_startofpacket),                      //                              .startofpacket
		.ff_rx_dval    (eth_tse_receive_valid),                              //                              .valid
		.ff_tx_data    (channel_adapter_0_out_data),                         //                      transmit.data
		.ff_tx_eop     (channel_adapter_0_out_endofpacket),                  //                              .endofpacket
		.ff_tx_err     (channel_adapter_0_out_error),                        //                              .error
		.ff_tx_mod     (channel_adapter_0_out_empty),                        //                              .empty
		.ff_tx_rdy     (channel_adapter_0_out_ready),                        //                              .ready
		.ff_tx_sop     (channel_adapter_0_out_startofpacket),                //                              .startofpacket
		.ff_tx_wren    (channel_adapter_0_out_valid),                        //                              .valid
		.mdc           (eth_tse_mac_mdio_connection_mdc),                    //           mac_mdio_connection.mdc
		.mdio_in       (eth_tse_mac_mdio_connection_mdio_in),                //                              .mdio_in
		.mdio_out      (eth_tse_mac_mdio_connection_mdio_out),               //                              .mdio_out
		.mdio_oen      (eth_tse_mac_mdio_connection_mdio_oen),               //                              .mdio_oen
		.magic_wakeup  (),                                                   //           mac_misc_connection.magic_wakeup
		.magic_sleep_n (),                                                   //                              .magic_sleep_n
		.ff_tx_crc_fwd (),                                                   //                              .ff_tx_crc_fwd
		.ff_tx_septy   (),                                                   //                              .ff_tx_septy
		.tx_ff_uflow   (),                                                   //                              .tx_ff_uflow
		.ff_tx_a_full  (),                                                   //                              .ff_tx_a_full
		.ff_tx_a_empty (),                                                   //                              .ff_tx_a_empty
		.rx_err_stat   (),                                                   //                              .rx_err_stat
		.rx_frm_type   (),                                                   //                              .rx_frm_type
		.ff_rx_dsav    (),                                                   //                              .ff_rx_dsav
		.ff_rx_a_full  (),                                                   //                              .ff_rx_a_full
		.ff_rx_a_empty ()                                                    //                              .ff_rx_a_empty
	);

	q_sys_ext_flash #(
		.DEVICE_FAMILY     ("MAX 10"),
		.CS_WIDTH          (1),
		.ADDR_WIDTH        (24),
		.ASI_WIDTH         (4),
		.ASMI_ADDR_WIDTH   (32),
		.ENABLE_4BYTE_ADDR (1),
		.IO_MODE           ("QUAD"),
		.CHIP_SELS         (1)
	) ext_flash (
		.clk                  (clock_bridge_0_in_clk_clk),                         //       clock_sink.clk
		.reset_n              (~rst_controller_005_reset_out_reset),               //            reset.reset_n
		.avl_csr_read         (mm_interconnect_1_ext_flash_avl_csr_read),          //          avl_csr.read
		.avl_csr_waitrequest  (mm_interconnect_1_ext_flash_avl_csr_waitrequest),   //                 .waitrequest
		.avl_csr_write        (mm_interconnect_1_ext_flash_avl_csr_write),         //                 .write
		.avl_csr_addr         (mm_interconnect_1_ext_flash_avl_csr_address),       //                 .address
		.avl_csr_wrdata       (mm_interconnect_1_ext_flash_avl_csr_writedata),     //                 .writedata
		.avl_csr_rddata       (mm_interconnect_1_ext_flash_avl_csr_readdata),      //                 .readdata
		.avl_csr_rddata_valid (mm_interconnect_1_ext_flash_avl_csr_readdatavalid), //                 .readdatavalid
		.avl_mem_write        (mm_interconnect_1_ext_flash_avl_mem_write),         //          avl_mem.write
		.avl_mem_burstcount   (mm_interconnect_1_ext_flash_avl_mem_burstcount),    //                 .burstcount
		.avl_mem_waitrequest  (mm_interconnect_1_ext_flash_avl_mem_waitrequest),   //                 .waitrequest
		.avl_mem_read         (mm_interconnect_1_ext_flash_avl_mem_read),          //                 .read
		.avl_mem_addr         (mm_interconnect_1_ext_flash_avl_mem_address),       //                 .address
		.avl_mem_wrdata       (mm_interconnect_1_ext_flash_avl_mem_writedata),     //                 .writedata
		.avl_mem_rddata       (mm_interconnect_1_ext_flash_avl_mem_readdata),      //                 .readdata
		.avl_mem_rddata_valid (mm_interconnect_1_ext_flash_avl_mem_readdatavalid), //                 .readdatavalid
		.avl_mem_byteenable   (mm_interconnect_1_ext_flash_avl_mem_byteenable),    //                 .byteenable
		.irq                  (irq_synchronizer_receiver_irq),                     // interrupt_sender.irq
		.flash_dataout        (ext_flash_flash_dataout_conduit_dataout),           //    flash_dataout.conduit_dataout
		.flash_dclk_out       (ext_flash_flash_dclk_out_conduit_dclk_out),         //   flash_dclk_out.conduit_dclk_out
		.flash_ncs            (ext_flash_flash_ncs_conduit_ncs)                    //        flash_ncs.conduit_ncs
	);

	q_sys_frame_timer frame_timer (
		.clk           (sys_clk_clk),                                 //           clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),         //         reset.reset_n
		.address       (mm_interconnect_1_frame_timer_s1_address),    //            s1.address
		.writedata     (mm_interconnect_1_frame_timer_s1_writedata),  //              .writedata
		.readdata      (mm_interconnect_1_frame_timer_s1_readdata),   //              .readdata
		.chipselect    (mm_interconnect_1_frame_timer_s1_chipselect), //              .chipselect
		.write_n       (~mm_interconnect_1_frame_timer_s1_write),     //              .write_n
		.irq           (),                                            //           irq.irq
		.timeout_pulse (frame_timer_export)                           // external_port.export
	);

	q_sys_msgdma_rx msgdma_rx (
		.mm_write_address                           (msgdma_rx_mm_write_address),                           //                mm_write.address
		.mm_write_write                             (msgdma_rx_mm_write_write),                             //                        .write
		.mm_write_byteenable                        (msgdma_rx_mm_write_byteenable),                        //                        .byteenable
		.mm_write_writedata                         (msgdma_rx_mm_write_writedata),                         //                        .writedata
		.mm_write_waitrequest                       (msgdma_rx_mm_write_waitrequest),                       //                        .waitrequest
		.descriptor_read_master_address             (msgdma_rx_descriptor_read_master_address),             //  descriptor_read_master.address
		.descriptor_read_master_read                (msgdma_rx_descriptor_read_master_read),                //                        .read
		.descriptor_read_master_readdata            (msgdma_rx_descriptor_read_master_readdata),            //                        .readdata
		.descriptor_read_master_waitrequest         (msgdma_rx_descriptor_read_master_waitrequest),         //                        .waitrequest
		.descriptor_read_master_readdatavalid       (msgdma_rx_descriptor_read_master_readdatavalid),       //                        .readdatavalid
		.descriptor_write_master_address            (msgdma_rx_descriptor_write_master_address),            // descriptor_write_master.address
		.descriptor_write_master_write              (msgdma_rx_descriptor_write_master_write),              //                        .write
		.descriptor_write_master_byteenable         (msgdma_rx_descriptor_write_master_byteenable),         //                        .byteenable
		.descriptor_write_master_writedata          (msgdma_rx_descriptor_write_master_writedata),          //                        .writedata
		.descriptor_write_master_waitrequest        (msgdma_rx_descriptor_write_master_waitrequest),        //                        .waitrequest
		.descriptor_write_master_response           (msgdma_rx_descriptor_write_master_response),           //                        .response
		.descriptor_write_master_writeresponsevalid (msgdma_rx_descriptor_write_master_writeresponsevalid), //                        .writeresponsevalid
		.clock_clk                                  (sys_clk_clk),                                          //                   clock.clk
		.reset_n_reset_n                            (~rst_controller_001_reset_out_reset),                  //                 reset_n.reset_n
		.csr_writedata                              (mm_interconnect_1_msgdma_rx_csr_writedata),            //                     csr.writedata
		.csr_write                                  (mm_interconnect_1_msgdma_rx_csr_write),                //                        .write
		.csr_byteenable                             (mm_interconnect_1_msgdma_rx_csr_byteenable),           //                        .byteenable
		.csr_readdata                               (mm_interconnect_1_msgdma_rx_csr_readdata),             //                        .readdata
		.csr_read                                   (mm_interconnect_1_msgdma_rx_csr_read),                 //                        .read
		.csr_address                                (mm_interconnect_1_msgdma_rx_csr_address),              //                        .address
		.prefetcher_csr_address                     (mm_interconnect_1_msgdma_rx_prefetcher_csr_address),   //          prefetcher_csr.address
		.prefetcher_csr_read                        (mm_interconnect_1_msgdma_rx_prefetcher_csr_read),      //                        .read
		.prefetcher_csr_write                       (mm_interconnect_1_msgdma_rx_prefetcher_csr_write),     //                        .write
		.prefetcher_csr_writedata                   (mm_interconnect_1_msgdma_rx_prefetcher_csr_writedata), //                        .writedata
		.prefetcher_csr_readdata                    (mm_interconnect_1_msgdma_rx_prefetcher_csr_readdata),  //                        .readdata
		.csr_irq_irq                                (irq_mapper_receiver1_irq),                             //                 csr_irq.irq
		.st_sink_data                               (avalon_st_adapter_001_out_0_data),                     //                 st_sink.data
		.st_sink_valid                              (avalon_st_adapter_001_out_0_valid),                    //                        .valid
		.st_sink_ready                              (avalon_st_adapter_001_out_0_ready),                    //                        .ready
		.st_sink_startofpacket                      (avalon_st_adapter_001_out_0_startofpacket),            //                        .startofpacket
		.st_sink_endofpacket                        (avalon_st_adapter_001_out_0_endofpacket),              //                        .endofpacket
		.st_sink_empty                              (avalon_st_adapter_001_out_0_empty),                    //                        .empty
		.st_sink_error                              (avalon_st_adapter_001_out_0_error)                     //                        .error
	);

	q_sys_msgdma_tx msgdma_tx (
		.mm_read_address                            (msgdma_tx_mm_read_address),                            //                 mm_read.address
		.mm_read_read                               (msgdma_tx_mm_read_read),                               //                        .read
		.mm_read_byteenable                         (msgdma_tx_mm_read_byteenable),                         //                        .byteenable
		.mm_read_readdata                           (msgdma_tx_mm_read_readdata),                           //                        .readdata
		.mm_read_waitrequest                        (msgdma_tx_mm_read_waitrequest),                        //                        .waitrequest
		.mm_read_readdatavalid                      (msgdma_tx_mm_read_readdatavalid),                      //                        .readdatavalid
		.descriptor_read_master_address             (msgdma_tx_descriptor_read_master_address),             //  descriptor_read_master.address
		.descriptor_read_master_read                (msgdma_tx_descriptor_read_master_read),                //                        .read
		.descriptor_read_master_readdata            (msgdma_tx_descriptor_read_master_readdata),            //                        .readdata
		.descriptor_read_master_waitrequest         (msgdma_tx_descriptor_read_master_waitrequest),         //                        .waitrequest
		.descriptor_read_master_readdatavalid       (msgdma_tx_descriptor_read_master_readdatavalid),       //                        .readdatavalid
		.descriptor_write_master_address            (msgdma_tx_descriptor_write_master_address),            // descriptor_write_master.address
		.descriptor_write_master_write              (msgdma_tx_descriptor_write_master_write),              //                        .write
		.descriptor_write_master_byteenable         (msgdma_tx_descriptor_write_master_byteenable),         //                        .byteenable
		.descriptor_write_master_writedata          (msgdma_tx_descriptor_write_master_writedata),          //                        .writedata
		.descriptor_write_master_waitrequest        (msgdma_tx_descriptor_write_master_waitrequest),        //                        .waitrequest
		.descriptor_write_master_response           (msgdma_tx_descriptor_write_master_response),           //                        .response
		.descriptor_write_master_writeresponsevalid (msgdma_tx_descriptor_write_master_writeresponsevalid), //                        .writeresponsevalid
		.clock_clk                                  (sys_clk_clk),                                          //                   clock.clk
		.reset_n_reset_n                            (~rst_controller_001_reset_out_reset),                  //                 reset_n.reset_n
		.csr_writedata                              (mm_interconnect_1_msgdma_tx_csr_writedata),            //                     csr.writedata
		.csr_write                                  (mm_interconnect_1_msgdma_tx_csr_write),                //                        .write
		.csr_byteenable                             (mm_interconnect_1_msgdma_tx_csr_byteenable),           //                        .byteenable
		.csr_readdata                               (mm_interconnect_1_msgdma_tx_csr_readdata),             //                        .readdata
		.csr_read                                   (mm_interconnect_1_msgdma_tx_csr_read),                 //                        .read
		.csr_address                                (mm_interconnect_1_msgdma_tx_csr_address),              //                        .address
		.prefetcher_csr_address                     (mm_interconnect_1_msgdma_tx_prefetcher_csr_address),   //          prefetcher_csr.address
		.prefetcher_csr_read                        (mm_interconnect_1_msgdma_tx_prefetcher_csr_read),      //                        .read
		.prefetcher_csr_write                       (mm_interconnect_1_msgdma_tx_prefetcher_csr_write),     //                        .write
		.prefetcher_csr_writedata                   (mm_interconnect_1_msgdma_tx_prefetcher_csr_writedata), //                        .writedata
		.prefetcher_csr_readdata                    (mm_interconnect_1_msgdma_tx_prefetcher_csr_readdata),  //                        .readdata
		.csr_irq_irq                                (irq_mapper_receiver0_irq),                             //                 csr_irq.irq
		.st_source_data                             (msgdma_tx_st_source_data),                             //               st_source.data
		.st_source_valid                            (msgdma_tx_st_source_valid),                            //                        .valid
		.st_source_ready                            (msgdma_tx_st_source_ready),                            //                        .ready
		.st_source_startofpacket                    (msgdma_tx_st_source_startofpacket),                    //                        .startofpacket
		.st_source_endofpacket                      (msgdma_tx_st_source_endofpacket),                      //                        .endofpacket
		.st_source_empty                            (msgdma_tx_st_source_empty),                            //                        .empty
		.st_source_error                            (msgdma_tx_st_source_error)                             //                        .error
	);

	altera_onchip_flash #(
		.INIT_FILENAME                       (""),
		.INIT_FILENAME_SIM                   (""),
		.DEVICE_FAMILY                       ("MAX 10"),
		.PART_NAME                           ("10M50DAF484C6GES"),
		.DEVICE_ID                           ("50"),
		.SECTOR1_START_ADDR                  (0),
		.SECTOR1_END_ADDR                    (8191),
		.SECTOR2_START_ADDR                  (8192),
		.SECTOR2_END_ADDR                    (16383),
		.SECTOR3_START_ADDR                  (16384),
		.SECTOR3_END_ADDR                    (114687),
		.SECTOR4_START_ADDR                  (114688),
		.SECTOR4_END_ADDR                    (188415),
		.SECTOR5_START_ADDR                  (188416),
		.SECTOR5_END_ADDR                    (360447),
		.MIN_VALID_ADDR                      (0),
		.MAX_VALID_ADDR                      (360447),
		.MIN_UFM_VALID_ADDR                  (0),
		.MAX_UFM_VALID_ADDR                  (114687),
		.SECTOR1_MAP                         (1),
		.SECTOR2_MAP                         (2),
		.SECTOR3_MAP                         (3),
		.SECTOR4_MAP                         (4),
		.SECTOR5_MAP                         (5),
		.ADDR_RANGE1_END_ADDR                (360447),
		.ADDR_RANGE2_END_ADDR                (360447),
		.ADDR_RANGE1_OFFSET                  (2048),
		.ADDR_RANGE2_OFFSET                  (0),
		.ADDR_RANGE3_OFFSET                  (0),
		.AVMM_DATA_ADDR_WIDTH                (19),
		.AVMM_DATA_DATA_WIDTH                (32),
		.AVMM_DATA_BURSTCOUNT_WIDTH          (4),
		.SECTOR_READ_PROTECTION_MODE         (0),
		.FLASH_SEQ_READ_DATA_COUNT           (4),
		.FLASH_ADDR_ALIGNMENT_BITS           (2),
		.FLASH_READ_CYCLE_MAX_INDEX          (5),
		.FLASH_RESET_CYCLE_MAX_INDEX         (12),
		.FLASH_BUSY_TIMEOUT_CYCLE_MAX_INDEX  (60),
		.FLASH_ERASE_TIMEOUT_CYCLE_MAX_INDEX (17500000),
		.FLASH_WRITE_TIMEOUT_CYCLE_MAX_INDEX (15250),
		.PARALLEL_MODE                       (1),
		.READ_AND_WRITE_MODE                 (1),
		.WRAPPING_BURST_MODE                 (0),
		.IS_DUAL_BOOT                        ("False"),
		.IS_ERAM_SKIP                        ("True"),
		.IS_COMPRESSED_IMAGE                 ("False")
	) onchip_flash (
		.clock                   (sys_clk_clk),                                       //    clk.clk
		.reset_n                 (~rst_controller_001_reset_out_reset),               // nreset.reset_n
		.avmm_data_addr          (mm_interconnect_1_onchip_flash_data_address),       //   data.address
		.avmm_data_read          (mm_interconnect_1_onchip_flash_data_read),          //       .read
		.avmm_data_writedata     (mm_interconnect_1_onchip_flash_data_writedata),     //       .writedata
		.avmm_data_write         (mm_interconnect_1_onchip_flash_data_write),         //       .write
		.avmm_data_readdata      (mm_interconnect_1_onchip_flash_data_readdata),      //       .readdata
		.avmm_data_waitrequest   (mm_interconnect_1_onchip_flash_data_waitrequest),   //       .waitrequest
		.avmm_data_readdatavalid (mm_interconnect_1_onchip_flash_data_readdatavalid), //       .readdatavalid
		.avmm_data_burstcount    (mm_interconnect_1_onchip_flash_data_burstcount),    //       .burstcount
		.avmm_csr_addr           (mm_interconnect_1_onchip_flash_csr_address),        //    csr.address
		.avmm_csr_read           (mm_interconnect_1_onchip_flash_csr_read),           //       .read
		.avmm_csr_writedata      (mm_interconnect_1_onchip_flash_csr_writedata),      //       .writedata
		.avmm_csr_write          (mm_interconnect_1_onchip_flash_csr_write),          //       .write
		.avmm_csr_readdata       (mm_interconnect_1_onchip_flash_csr_readdata)        //       .readdata
	);

	q_sys_output_pio output_pio (
		.clk        (sys_clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_004_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_1_output_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_output_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_output_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_output_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_output_pio_s1_readdata),   //                    .readdata
		.out_port   (led_pio_external_connection_export)          // external_connection.export
	);

	sensor_algo sensor_interface (
		.csr_address            (mm_interconnect_1_sensor_interface_csr_address),         //                       csr.address
		.csr_read               (mm_interconnect_1_sensor_interface_csr_read),            //                          .read
		.csr_readdata           (mm_interconnect_1_sensor_interface_csr_readdata),        //                          .readdata
		.csr_write              (mm_interconnect_1_sensor_interface_csr_write),           //                          .write
		.csr_writedata          (mm_interconnect_1_sensor_interface_csr_writedata),       //                          .writedata
		.csr_byteenable         (mm_interconnect_1_sensor_interface_csr_byteenable),      //                          .byteenable
		.data_out_endofpacket   (sensor_interface_data_out_endofpacket),                  //                  data_out.endofpacket
		.data_out_data          (sensor_interface_data_out_data),                         //                          .data
		.data_out_empty         (sensor_interface_data_out_empty),                        //                          .empty
		.data_out_ready         (sensor_interface_data_out_ready),                        //                          .ready
		.data_out_startofpacket (sensor_interface_data_out_startofpacket),                //                          .startofpacket
		.data_out_valid         (sensor_interface_data_out_valid),                        //                          .valid
		.clk_clk                (sys_clk_clk),                                            //                       clk.clk
		.rst_reset              (rst_controller_001_reset_out_reset),                     //                       rst.reset
		.in_adc_data            (sensor_in_adc_data),                                     //                    sensor.in_adc_data
		.in_trg                 (sensor_in_trg),                                          //                          .in_trg
		.out_adc_clk            (sensor_out_adc_clk),                                     //                          .out_adc_clk
		.out_adc_cnv            (sensor_out_adc_cnv),                                     //                          .out_adc_cnv
		.out_sensor_clk         (sensor_out_sensor_clk),                                  //                          .out_sensor_clk
		.out_sensor_gain        (sensor_out_sensor_gain),                                 //                          .out_sensor_gain
		.out_sensor_rst         (sensor_out_sensor_rst),                                  //                          .out_sensor_rst
		.status_out             (sensor_status_status_out),                               //                status_out.status_out
		.ext_input              (sensor_synchro_ext_input),                               //                   synchro.ext_input
		.serial_rx              (sensor_synchro_serial_rx),                               //                          .serial_rx
		.serial_tx              (sensor_synchro_serial_tx),                               //                          .serial_tx
		.address                (sensor_interface_calibration_ram_interface_address),     // calibration_ram_interface.address
		.clken                  (sensor_interface_calibration_ram_interface_read),        //                          .read
		.cali_fac               (sensor_interface_calibration_ram_interface_readdata),    //                          .readdata
		.waitrequest            (sensor_interface_calibration_ram_interface_waitrequest)  //                          .waitrequest
	);

	q_sys_sys_clk_timer sys_clk_timer (
		.clk        (sys_clk_clk),                                   //   clk.clk
		.reset_n    (~rst_controller_004_reset_out_reset),           // reset.reset_n
		.address    (mm_interconnect_1_sys_clk_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_sys_clk_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_sys_clk_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_sys_clk_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_sys_clk_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                       //   irq.irq
	);

	q_sys_sysid sysid (
		.clock    (sys_clk_clk),                                    //           clk.clk
		.reset_n  (~rst_controller_004_reset_out_reset),            //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_control_slave_address)   //              .address
	);

	q_sys_tx_multiplexer tx_multiplexer (
		.clk               (sys_clk_clk),                           //   clk.clk
		.reset_n           (~rst_controller_001_reset_out_reset),   // reset.reset_n
		.out_data          (tx_multiplexer_out_data),               //   out.data
		.out_valid         (tx_multiplexer_out_valid),              //      .valid
		.out_ready         (tx_multiplexer_out_ready),              //      .ready
		.out_startofpacket (tx_multiplexer_out_startofpacket),      //      .startofpacket
		.out_endofpacket   (tx_multiplexer_out_endofpacket),        //      .endofpacket
		.out_empty         (tx_multiplexer_out_empty),              //      .empty
		.out_error         (tx_multiplexer_out_error),              //      .error
		.out_channel       (tx_multiplexer_out_channel),            //      .channel
		.in0_data          (msgdma_tx_st_source_data),              //   in0.data
		.in0_valid         (msgdma_tx_st_source_valid),             //      .valid
		.in0_ready         (msgdma_tx_st_source_ready),             //      .ready
		.in0_startofpacket (msgdma_tx_st_source_startofpacket),     //      .startofpacket
		.in0_endofpacket   (msgdma_tx_st_source_endofpacket),       //      .endofpacket
		.in0_empty         (msgdma_tx_st_source_empty),             //      .empty
		.in0_error         (msgdma_tx_st_source_error),             //      .error
		.in1_data          (avalon_st_adapter_out_0_data),          //   in1.data
		.in1_valid         (avalon_st_adapter_out_0_valid),         //      .valid
		.in1_ready         (avalon_st_adapter_out_0_ready),         //      .ready
		.in1_startofpacket (avalon_st_adapter_out_0_startofpacket), //      .startofpacket
		.in1_endofpacket   (avalon_st_adapter_out_0_endofpacket),   //      .endofpacket
		.in1_empty         (avalon_st_adapter_out_0_empty),         //      .empty
		.in1_error         (avalon_st_adapter_out_0_error)          //      .error
	);

	udp_generator udp_generator (
		.clk_clk                (sys_clk_clk),                                    //      clk.clk
		.rst_reset              (rst_controller_001_reset_out_reset),             //      rst.reset
		.csr_address            (mm_interconnect_1_udp_generator_csr_address),    //      csr.address
		.csr_write              (mm_interconnect_1_udp_generator_csr_write),      //         .write
		.csr_writedata          (mm_interconnect_1_udp_generator_csr_writedata),  //         .writedata
		.csr_byteenable         (mm_interconnect_1_udp_generator_csr_byteenable), //         .byteenable
		.csr_read               (mm_interconnect_1_udp_generator_csr_read),       //         .read
		.csr_readdata           (mm_interconnect_1_udp_generator_csr_readdata),   //         .readdata
		.data_in_data           (sensor_interface_data_out_data),                 //  data_in.data
		.data_in_ready          (sensor_interface_data_out_ready),                //         .ready
		.data_in_valid          (sensor_interface_data_out_valid),                //         .valid
		.data_in_empty          (sensor_interface_data_out_empty),                //         .empty
		.data_in_endofpacket    (sensor_interface_data_out_endofpacket),          //         .endofpacket
		.data_in_startofpacket  (sensor_interface_data_out_startofpacket),        //         .startofpacket
		.data_out_data          (udp_generator_data_out_data),                    // data_out.data
		.data_out_empty         (udp_generator_data_out_empty),                   //         .empty
		.data_out_endofpacket   (udp_generator_data_out_endofpacket),             //         .endofpacket
		.data_out_startofpacket (udp_generator_data_out_startofpacket),           //         .startofpacket
		.data_out_ready         (udp_generator_data_out_ready),                   //         .ready
		.data_out_valid         (udp_generator_data_out_valid)                    //         .valid
	);

	q_sys_mm_interconnect_0 mm_interconnect_0 (
		.sys_clk_clk_clk                                        (sys_clk_clk),                                            //                                sys_clk_clk.clk
		.sensor_interface_rst_reset_bridge_in_reset_reset       (rst_controller_001_reset_out_reset),                     // sensor_interface_rst_reset_bridge_in_reset.reset
		.sensor_interface_calibration_ram_interface_address     (sensor_interface_calibration_ram_interface_address),     // sensor_interface_calibration_ram_interface.address
		.sensor_interface_calibration_ram_interface_waitrequest (sensor_interface_calibration_ram_interface_waitrequest), //                                           .waitrequest
		.sensor_interface_calibration_ram_interface_read        (sensor_interface_calibration_ram_interface_read),        //                                           .read
		.sensor_interface_calibration_ram_interface_readdata    (sensor_interface_calibration_ram_interface_readdata),    //                                           .readdata
		.calibration_ram_s2_address                             (mm_interconnect_0_calibration_ram_s2_address),           //                         calibration_ram_s2.address
		.calibration_ram_s2_write                               (mm_interconnect_0_calibration_ram_s2_write),             //                                           .write
		.calibration_ram_s2_readdata                            (mm_interconnect_0_calibration_ram_s2_readdata),          //                                           .readdata
		.calibration_ram_s2_writedata                           (mm_interconnect_0_calibration_ram_s2_writedata),         //                                           .writedata
		.calibration_ram_s2_byteenable                          (mm_interconnect_0_calibration_ram_s2_byteenable),        //                                           .byteenable
		.calibration_ram_s2_chipselect                          (mm_interconnect_0_calibration_ram_s2_chipselect),        //                                           .chipselect
		.calibration_ram_s2_clken                               (mm_interconnect_0_calibration_ram_s2_clken)              //                                           .clken
	);

	q_sys_mm_interconnect_1 mm_interconnect_1 (
		.ddr3_ram_afi_clk_clk                                      (ddr3_ram_afi_clk_clk),                                 //                                    ddr3_ram_afi_clk.clk
		.ext_flash_clock_bridge_out_clk_clk                        (clock_bridge_0_in_clk_clk),                            //                      ext_flash_clock_bridge_out_clk.clk
		.sys_clk_clk_clk                                           (sys_clk_clk),                                          //                                         sys_clk_clk.clk
		.cpu_reset_reset_bridge_in_reset_reset                     (rst_controller_001_reset_out_reset),                   //                     cpu_reset_reset_bridge_in_reset.reset
		.ddr3_ram_avl_translator_reset_reset_bridge_in_reset_reset (rst_controller_006_reset_out_reset),                   // ddr3_ram_avl_translator_reset_reset_bridge_in_reset.reset
		.ddr3_ram_soft_reset_reset_bridge_in_reset_reset           (rst_controller_006_reset_out_reset),                   //           ddr3_ram_soft_reset_reset_bridge_in_reset.reset
		.eth_tse_reset_connection_reset_bridge_in_reset_reset      (rst_controller_004_reset_out_reset),                   //      eth_tse_reset_connection_reset_bridge_in_reset.reset
		.ext_flash_reset_reset_bridge_in_reset_reset               (rst_controller_005_reset_out_reset),                   //               ext_flash_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                                   (cpu_data_master_address),                              //                                     cpu_data_master.address
		.cpu_data_master_waitrequest                               (cpu_data_master_waitrequest),                          //                                                    .waitrequest
		.cpu_data_master_byteenable                                (cpu_data_master_byteenable),                           //                                                    .byteenable
		.cpu_data_master_read                                      (cpu_data_master_read),                                 //                                                    .read
		.cpu_data_master_readdata                                  (cpu_data_master_readdata),                             //                                                    .readdata
		.cpu_data_master_readdatavalid                             (cpu_data_master_readdatavalid),                        //                                                    .readdatavalid
		.cpu_data_master_write                                     (cpu_data_master_write),                                //                                                    .write
		.cpu_data_master_writedata                                 (cpu_data_master_writedata),                            //                                                    .writedata
		.cpu_data_master_debugaccess                               (cpu_data_master_debugaccess),                          //                                                    .debugaccess
		.cpu_instruction_master_address                            (cpu_instruction_master_address),                       //                              cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                        (cpu_instruction_master_waitrequest),                   //                                                    .waitrequest
		.cpu_instruction_master_read                               (cpu_instruction_master_read),                          //                                                    .read
		.cpu_instruction_master_readdata                           (cpu_instruction_master_readdata),                      //                                                    .readdata
		.cpu_instruction_master_readdatavalid                      (cpu_instruction_master_readdatavalid),                 //                                                    .readdatavalid
		.msgdma_rx_descriptor_read_master_address                  (msgdma_rx_descriptor_read_master_address),             //                    msgdma_rx_descriptor_read_master.address
		.msgdma_rx_descriptor_read_master_waitrequest              (msgdma_rx_descriptor_read_master_waitrequest),         //                                                    .waitrequest
		.msgdma_rx_descriptor_read_master_read                     (msgdma_rx_descriptor_read_master_read),                //                                                    .read
		.msgdma_rx_descriptor_read_master_readdata                 (msgdma_rx_descriptor_read_master_readdata),            //                                                    .readdata
		.msgdma_rx_descriptor_read_master_readdatavalid            (msgdma_rx_descriptor_read_master_readdatavalid),       //                                                    .readdatavalid
		.msgdma_rx_descriptor_write_master_address                 (msgdma_rx_descriptor_write_master_address),            //                   msgdma_rx_descriptor_write_master.address
		.msgdma_rx_descriptor_write_master_waitrequest             (msgdma_rx_descriptor_write_master_waitrequest),        //                                                    .waitrequest
		.msgdma_rx_descriptor_write_master_byteenable              (msgdma_rx_descriptor_write_master_byteenable),         //                                                    .byteenable
		.msgdma_rx_descriptor_write_master_write                   (msgdma_rx_descriptor_write_master_write),              //                                                    .write
		.msgdma_rx_descriptor_write_master_writedata               (msgdma_rx_descriptor_write_master_writedata),          //                                                    .writedata
		.msgdma_rx_descriptor_write_master_response                (msgdma_rx_descriptor_write_master_response),           //                                                    .response
		.msgdma_rx_descriptor_write_master_writeresponsevalid      (msgdma_rx_descriptor_write_master_writeresponsevalid), //                                                    .writeresponsevalid
		.msgdma_rx_mm_write_address                                (msgdma_rx_mm_write_address),                           //                                  msgdma_rx_mm_write.address
		.msgdma_rx_mm_write_waitrequest                            (msgdma_rx_mm_write_waitrequest),                       //                                                    .waitrequest
		.msgdma_rx_mm_write_byteenable                             (msgdma_rx_mm_write_byteenable),                        //                                                    .byteenable
		.msgdma_rx_mm_write_write                                  (msgdma_rx_mm_write_write),                             //                                                    .write
		.msgdma_rx_mm_write_writedata                              (msgdma_rx_mm_write_writedata),                         //                                                    .writedata
		.msgdma_tx_descriptor_read_master_address                  (msgdma_tx_descriptor_read_master_address),             //                    msgdma_tx_descriptor_read_master.address
		.msgdma_tx_descriptor_read_master_waitrequest              (msgdma_tx_descriptor_read_master_waitrequest),         //                                                    .waitrequest
		.msgdma_tx_descriptor_read_master_read                     (msgdma_tx_descriptor_read_master_read),                //                                                    .read
		.msgdma_tx_descriptor_read_master_readdata                 (msgdma_tx_descriptor_read_master_readdata),            //                                                    .readdata
		.msgdma_tx_descriptor_read_master_readdatavalid            (msgdma_tx_descriptor_read_master_readdatavalid),       //                                                    .readdatavalid
		.msgdma_tx_descriptor_write_master_address                 (msgdma_tx_descriptor_write_master_address),            //                   msgdma_tx_descriptor_write_master.address
		.msgdma_tx_descriptor_write_master_waitrequest             (msgdma_tx_descriptor_write_master_waitrequest),        //                                                    .waitrequest
		.msgdma_tx_descriptor_write_master_byteenable              (msgdma_tx_descriptor_write_master_byteenable),         //                                                    .byteenable
		.msgdma_tx_descriptor_write_master_write                   (msgdma_tx_descriptor_write_master_write),              //                                                    .write
		.msgdma_tx_descriptor_write_master_writedata               (msgdma_tx_descriptor_write_master_writedata),          //                                                    .writedata
		.msgdma_tx_descriptor_write_master_response                (msgdma_tx_descriptor_write_master_response),           //                                                    .response
		.msgdma_tx_descriptor_write_master_writeresponsevalid      (msgdma_tx_descriptor_write_master_writeresponsevalid), //                                                    .writeresponsevalid
		.msgdma_tx_mm_read_address                                 (msgdma_tx_mm_read_address),                            //                                   msgdma_tx_mm_read.address
		.msgdma_tx_mm_read_waitrequest                             (msgdma_tx_mm_read_waitrequest),                        //                                                    .waitrequest
		.msgdma_tx_mm_read_byteenable                              (msgdma_tx_mm_read_byteenable),                         //                                                    .byteenable
		.msgdma_tx_mm_read_read                                    (msgdma_tx_mm_read_read),                               //                                                    .read
		.msgdma_tx_mm_read_readdata                                (msgdma_tx_mm_read_readdata),                           //                                                    .readdata
		.msgdma_tx_mm_read_readdatavalid                           (msgdma_tx_mm_read_readdatavalid),                      //                                                    .readdatavalid
		.button_pio_s1_address                                     (mm_interconnect_1_button_pio_s1_address),              //                                       button_pio_s1.address
		.button_pio_s1_readdata                                    (mm_interconnect_1_button_pio_s1_readdata),             //                                                    .readdata
		.calibration_ram_s1_address                                (mm_interconnect_1_calibration_ram_s1_address),         //                                  calibration_ram_s1.address
		.calibration_ram_s1_write                                  (mm_interconnect_1_calibration_ram_s1_write),           //                                                    .write
		.calibration_ram_s1_readdata                               (mm_interconnect_1_calibration_ram_s1_readdata),        //                                                    .readdata
		.calibration_ram_s1_writedata                              (mm_interconnect_1_calibration_ram_s1_writedata),       //                                                    .writedata
		.calibration_ram_s1_byteenable                             (mm_interconnect_1_calibration_ram_s1_byteenable),      //                                                    .byteenable
		.calibration_ram_s1_chipselect                             (mm_interconnect_1_calibration_ram_s1_chipselect),      //                                                    .chipselect
		.calibration_ram_s1_clken                                  (mm_interconnect_1_calibration_ram_s1_clken),           //                                                    .clken
		.cpu_debug_mem_slave_address                               (mm_interconnect_1_cpu_debug_mem_slave_address),        //                                 cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write                                 (mm_interconnect_1_cpu_debug_mem_slave_write),          //                                                    .write
		.cpu_debug_mem_slave_read                                  (mm_interconnect_1_cpu_debug_mem_slave_read),           //                                                    .read
		.cpu_debug_mem_slave_readdata                              (mm_interconnect_1_cpu_debug_mem_slave_readdata),       //                                                    .readdata
		.cpu_debug_mem_slave_writedata                             (mm_interconnect_1_cpu_debug_mem_slave_writedata),      //                                                    .writedata
		.cpu_debug_mem_slave_byteenable                            (mm_interconnect_1_cpu_debug_mem_slave_byteenable),     //                                                    .byteenable
		.cpu_debug_mem_slave_waitrequest                           (mm_interconnect_1_cpu_debug_mem_slave_waitrequest),    //                                                    .waitrequest
		.cpu_debug_mem_slave_debugaccess                           (mm_interconnect_1_cpu_debug_mem_slave_debugaccess),    //                                                    .debugaccess
		.ddr3_ram_avl_address                                      (mm_interconnect_1_ddr3_ram_avl_address),               //                                        ddr3_ram_avl.address
		.ddr3_ram_avl_write                                        (mm_interconnect_1_ddr3_ram_avl_write),                 //                                                    .write
		.ddr3_ram_avl_read                                         (mm_interconnect_1_ddr3_ram_avl_read),                  //                                                    .read
		.ddr3_ram_avl_readdata                                     (mm_interconnect_1_ddr3_ram_avl_readdata),              //                                                    .readdata
		.ddr3_ram_avl_writedata                                    (mm_interconnect_1_ddr3_ram_avl_writedata),             //                                                    .writedata
		.ddr3_ram_avl_beginbursttransfer                           (mm_interconnect_1_ddr3_ram_avl_beginbursttransfer),    //                                                    .beginbursttransfer
		.ddr3_ram_avl_burstcount                                   (mm_interconnect_1_ddr3_ram_avl_burstcount),            //                                                    .burstcount
		.ddr3_ram_avl_byteenable                                   (mm_interconnect_1_ddr3_ram_avl_byteenable),            //                                                    .byteenable
		.ddr3_ram_avl_readdatavalid                                (mm_interconnect_1_ddr3_ram_avl_readdatavalid),         //                                                    .readdatavalid
		.ddr3_ram_avl_waitrequest                                  (~mm_interconnect_1_ddr3_ram_avl_waitrequest),          //                                                    .waitrequest
		.debug_uart_s1_address                                     (mm_interconnect_1_debug_uart_s1_address),              //                                       debug_uart_s1.address
		.debug_uart_s1_write                                       (mm_interconnect_1_debug_uart_s1_write),                //                                                    .write
		.debug_uart_s1_read                                        (mm_interconnect_1_debug_uart_s1_read),                 //                                                    .read
		.debug_uart_s1_readdata                                    (mm_interconnect_1_debug_uart_s1_readdata),             //                                                    .readdata
		.debug_uart_s1_writedata                                   (mm_interconnect_1_debug_uart_s1_writedata),            //                                                    .writedata
		.debug_uart_s1_begintransfer                               (mm_interconnect_1_debug_uart_s1_begintransfer),        //                                                    .begintransfer
		.debug_uart_s1_chipselect                                  (mm_interconnect_1_debug_uart_s1_chipselect),           //                                                    .chipselect
		.descriptor_memory_s1_address                              (mm_interconnect_1_descriptor_memory_s1_address),       //                                descriptor_memory_s1.address
		.descriptor_memory_s1_write                                (mm_interconnect_1_descriptor_memory_s1_write),         //                                                    .write
		.descriptor_memory_s1_readdata                             (mm_interconnect_1_descriptor_memory_s1_readdata),      //                                                    .readdata
		.descriptor_memory_s1_writedata                            (mm_interconnect_1_descriptor_memory_s1_writedata),     //                                                    .writedata
		.descriptor_memory_s1_byteenable                           (mm_interconnect_1_descriptor_memory_s1_byteenable),    //                                                    .byteenable
		.descriptor_memory_s1_chipselect                           (mm_interconnect_1_descriptor_memory_s1_chipselect),    //                                                    .chipselect
		.descriptor_memory_s1_clken                                (mm_interconnect_1_descriptor_memory_s1_clken),         //                                                    .clken
		.eth_tse_control_port_address                              (mm_interconnect_1_eth_tse_control_port_address),       //                                eth_tse_control_port.address
		.eth_tse_control_port_write                                (mm_interconnect_1_eth_tse_control_port_write),         //                                                    .write
		.eth_tse_control_port_read                                 (mm_interconnect_1_eth_tse_control_port_read),          //                                                    .read
		.eth_tse_control_port_readdata                             (mm_interconnect_1_eth_tse_control_port_readdata),      //                                                    .readdata
		.eth_tse_control_port_writedata                            (mm_interconnect_1_eth_tse_control_port_writedata),     //                                                    .writedata
		.eth_tse_control_port_waitrequest                          (mm_interconnect_1_eth_tse_control_port_waitrequest),   //                                                    .waitrequest
		.ext_flash_avl_csr_address                                 (mm_interconnect_1_ext_flash_avl_csr_address),          //                                   ext_flash_avl_csr.address
		.ext_flash_avl_csr_write                                   (mm_interconnect_1_ext_flash_avl_csr_write),            //                                                    .write
		.ext_flash_avl_csr_read                                    (mm_interconnect_1_ext_flash_avl_csr_read),             //                                                    .read
		.ext_flash_avl_csr_readdata                                (mm_interconnect_1_ext_flash_avl_csr_readdata),         //                                                    .readdata
		.ext_flash_avl_csr_writedata                               (mm_interconnect_1_ext_flash_avl_csr_writedata),        //                                                    .writedata
		.ext_flash_avl_csr_readdatavalid                           (mm_interconnect_1_ext_flash_avl_csr_readdatavalid),    //                                                    .readdatavalid
		.ext_flash_avl_csr_waitrequest                             (mm_interconnect_1_ext_flash_avl_csr_waitrequest),      //                                                    .waitrequest
		.ext_flash_avl_mem_address                                 (mm_interconnect_1_ext_flash_avl_mem_address),          //                                   ext_flash_avl_mem.address
		.ext_flash_avl_mem_write                                   (mm_interconnect_1_ext_flash_avl_mem_write),            //                                                    .write
		.ext_flash_avl_mem_read                                    (mm_interconnect_1_ext_flash_avl_mem_read),             //                                                    .read
		.ext_flash_avl_mem_readdata                                (mm_interconnect_1_ext_flash_avl_mem_readdata),         //                                                    .readdata
		.ext_flash_avl_mem_writedata                               (mm_interconnect_1_ext_flash_avl_mem_writedata),        //                                                    .writedata
		.ext_flash_avl_mem_burstcount                              (mm_interconnect_1_ext_flash_avl_mem_burstcount),       //                                                    .burstcount
		.ext_flash_avl_mem_byteenable                              (mm_interconnect_1_ext_flash_avl_mem_byteenable),       //                                                    .byteenable
		.ext_flash_avl_mem_readdatavalid                           (mm_interconnect_1_ext_flash_avl_mem_readdatavalid),    //                                                    .readdatavalid
		.ext_flash_avl_mem_waitrequest                             (mm_interconnect_1_ext_flash_avl_mem_waitrequest),      //                                                    .waitrequest
		.frame_timer_s1_address                                    (mm_interconnect_1_frame_timer_s1_address),             //                                      frame_timer_s1.address
		.frame_timer_s1_write                                      (mm_interconnect_1_frame_timer_s1_write),               //                                                    .write
		.frame_timer_s1_readdata                                   (mm_interconnect_1_frame_timer_s1_readdata),            //                                                    .readdata
		.frame_timer_s1_writedata                                  (mm_interconnect_1_frame_timer_s1_writedata),           //                                                    .writedata
		.frame_timer_s1_chipselect                                 (mm_interconnect_1_frame_timer_s1_chipselect),          //                                                    .chipselect
		.msgdma_rx_csr_address                                     (mm_interconnect_1_msgdma_rx_csr_address),              //                                       msgdma_rx_csr.address
		.msgdma_rx_csr_write                                       (mm_interconnect_1_msgdma_rx_csr_write),                //                                                    .write
		.msgdma_rx_csr_read                                        (mm_interconnect_1_msgdma_rx_csr_read),                 //                                                    .read
		.msgdma_rx_csr_readdata                                    (mm_interconnect_1_msgdma_rx_csr_readdata),             //                                                    .readdata
		.msgdma_rx_csr_writedata                                   (mm_interconnect_1_msgdma_rx_csr_writedata),            //                                                    .writedata
		.msgdma_rx_csr_byteenable                                  (mm_interconnect_1_msgdma_rx_csr_byteenable),           //                                                    .byteenable
		.msgdma_rx_prefetcher_csr_address                          (mm_interconnect_1_msgdma_rx_prefetcher_csr_address),   //                            msgdma_rx_prefetcher_csr.address
		.msgdma_rx_prefetcher_csr_write                            (mm_interconnect_1_msgdma_rx_prefetcher_csr_write),     //                                                    .write
		.msgdma_rx_prefetcher_csr_read                             (mm_interconnect_1_msgdma_rx_prefetcher_csr_read),      //                                                    .read
		.msgdma_rx_prefetcher_csr_readdata                         (mm_interconnect_1_msgdma_rx_prefetcher_csr_readdata),  //                                                    .readdata
		.msgdma_rx_prefetcher_csr_writedata                        (mm_interconnect_1_msgdma_rx_prefetcher_csr_writedata), //                                                    .writedata
		.msgdma_tx_csr_address                                     (mm_interconnect_1_msgdma_tx_csr_address),              //                                       msgdma_tx_csr.address
		.msgdma_tx_csr_write                                       (mm_interconnect_1_msgdma_tx_csr_write),                //                                                    .write
		.msgdma_tx_csr_read                                        (mm_interconnect_1_msgdma_tx_csr_read),                 //                                                    .read
		.msgdma_tx_csr_readdata                                    (mm_interconnect_1_msgdma_tx_csr_readdata),             //                                                    .readdata
		.msgdma_tx_csr_writedata                                   (mm_interconnect_1_msgdma_tx_csr_writedata),            //                                                    .writedata
		.msgdma_tx_csr_byteenable                                  (mm_interconnect_1_msgdma_tx_csr_byteenable),           //                                                    .byteenable
		.msgdma_tx_prefetcher_csr_address                          (mm_interconnect_1_msgdma_tx_prefetcher_csr_address),   //                            msgdma_tx_prefetcher_csr.address
		.msgdma_tx_prefetcher_csr_write                            (mm_interconnect_1_msgdma_tx_prefetcher_csr_write),     //                                                    .write
		.msgdma_tx_prefetcher_csr_read                             (mm_interconnect_1_msgdma_tx_prefetcher_csr_read),      //                                                    .read
		.msgdma_tx_prefetcher_csr_readdata                         (mm_interconnect_1_msgdma_tx_prefetcher_csr_readdata),  //                                                    .readdata
		.msgdma_tx_prefetcher_csr_writedata                        (mm_interconnect_1_msgdma_tx_prefetcher_csr_writedata), //                                                    .writedata
		.onchip_flash_csr_address                                  (mm_interconnect_1_onchip_flash_csr_address),           //                                    onchip_flash_csr.address
		.onchip_flash_csr_write                                    (mm_interconnect_1_onchip_flash_csr_write),             //                                                    .write
		.onchip_flash_csr_read                                     (mm_interconnect_1_onchip_flash_csr_read),              //                                                    .read
		.onchip_flash_csr_readdata                                 (mm_interconnect_1_onchip_flash_csr_readdata),          //                                                    .readdata
		.onchip_flash_csr_writedata                                (mm_interconnect_1_onchip_flash_csr_writedata),         //                                                    .writedata
		.onchip_flash_data_address                                 (mm_interconnect_1_onchip_flash_data_address),          //                                   onchip_flash_data.address
		.onchip_flash_data_write                                   (mm_interconnect_1_onchip_flash_data_write),            //                                                    .write
		.onchip_flash_data_read                                    (mm_interconnect_1_onchip_flash_data_read),             //                                                    .read
		.onchip_flash_data_readdata                                (mm_interconnect_1_onchip_flash_data_readdata),         //                                                    .readdata
		.onchip_flash_data_writedata                               (mm_interconnect_1_onchip_flash_data_writedata),        //                                                    .writedata
		.onchip_flash_data_burstcount                              (mm_interconnect_1_onchip_flash_data_burstcount),       //                                                    .burstcount
		.onchip_flash_data_readdatavalid                           (mm_interconnect_1_onchip_flash_data_readdatavalid),    //                                                    .readdatavalid
		.onchip_flash_data_waitrequest                             (mm_interconnect_1_onchip_flash_data_waitrequest),      //                                                    .waitrequest
		.output_pio_s1_address                                     (mm_interconnect_1_output_pio_s1_address),              //                                       output_pio_s1.address
		.output_pio_s1_write                                       (mm_interconnect_1_output_pio_s1_write),                //                                                    .write
		.output_pio_s1_readdata                                    (mm_interconnect_1_output_pio_s1_readdata),             //                                                    .readdata
		.output_pio_s1_writedata                                   (mm_interconnect_1_output_pio_s1_writedata),            //                                                    .writedata
		.output_pio_s1_chipselect                                  (mm_interconnect_1_output_pio_s1_chipselect),           //                                                    .chipselect
		.sensor_interface_csr_address                              (mm_interconnect_1_sensor_interface_csr_address),       //                                sensor_interface_csr.address
		.sensor_interface_csr_write                                (mm_interconnect_1_sensor_interface_csr_write),         //                                                    .write
		.sensor_interface_csr_read                                 (mm_interconnect_1_sensor_interface_csr_read),          //                                                    .read
		.sensor_interface_csr_readdata                             (mm_interconnect_1_sensor_interface_csr_readdata),      //                                                    .readdata
		.sensor_interface_csr_writedata                            (mm_interconnect_1_sensor_interface_csr_writedata),     //                                                    .writedata
		.sensor_interface_csr_byteenable                           (mm_interconnect_1_sensor_interface_csr_byteenable),    //                                                    .byteenable
		.sys_clk_timer_s1_address                                  (mm_interconnect_1_sys_clk_timer_s1_address),           //                                    sys_clk_timer_s1.address
		.sys_clk_timer_s1_write                                    (mm_interconnect_1_sys_clk_timer_s1_write),             //                                                    .write
		.sys_clk_timer_s1_readdata                                 (mm_interconnect_1_sys_clk_timer_s1_readdata),          //                                                    .readdata
		.sys_clk_timer_s1_writedata                                (mm_interconnect_1_sys_clk_timer_s1_writedata),         //                                                    .writedata
		.sys_clk_timer_s1_chipselect                               (mm_interconnect_1_sys_clk_timer_s1_chipselect),        //                                                    .chipselect
		.sysid_control_slave_address                               (mm_interconnect_1_sysid_control_slave_address),        //                                 sysid_control_slave.address
		.sysid_control_slave_readdata                              (mm_interconnect_1_sysid_control_slave_readdata),       //                                                    .readdata
		.udp_generator_csr_address                                 (mm_interconnect_1_udp_generator_csr_address),          //                                   udp_generator_csr.address
		.udp_generator_csr_write                                   (mm_interconnect_1_udp_generator_csr_write),            //                                                    .write
		.udp_generator_csr_read                                    (mm_interconnect_1_udp_generator_csr_read),             //                                                    .read
		.udp_generator_csr_readdata                                (mm_interconnect_1_udp_generator_csr_readdata),         //                                                    .readdata
		.udp_generator_csr_writedata                               (mm_interconnect_1_udp_generator_csr_writedata),        //                                                    .writedata
		.udp_generator_csr_byteenable                              (mm_interconnect_1_udp_generator_csr_byteenable)        //                                                    .byteenable
	);

	q_sys_irq_mapper irq_mapper (
		.clk           (sys_clk_clk),                        //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.sender_irq    (cpu_irq_irq)                         //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (clock_bridge_0_in_clk_clk),          //       receiver_clk.clk
		.sender_clk     (sys_clk_clk),                        //         sender_clk.clk
		.receiver_reset (rst_controller_005_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	q_sys_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (1),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (sys_clk_clk),                           // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_001_reset_out_reset),    // in_rst_0.reset
		.in_0_data           (udp_generator_data_out_data),           //     in_0.data
		.in_0_valid          (udp_generator_data_out_valid),          //         .valid
		.in_0_ready          (udp_generator_data_out_ready),          //         .ready
		.in_0_startofpacket  (udp_generator_data_out_startofpacket),  //         .startofpacket
		.in_0_endofpacket    (udp_generator_data_out_endofpacket),    //         .endofpacket
		.in_0_empty          (udp_generator_data_out_empty),          //         .empty
		.out_0_data          (avalon_st_adapter_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_out_0_empty),         //         .empty
		.out_0_error         (avalon_st_adapter_out_0_error)          //         .error
	);

	q_sys_avalon_st_adapter_001 #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (6),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (2),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (6),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_001 (
		.in_clk_0_clk        (sys_clk_clk),                               // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_004_reset_out_reset),        // in_rst_0.reset
		.in_0_data           (eth_tse_receive_data),                      //     in_0.data
		.in_0_valid          (eth_tse_receive_valid),                     //         .valid
		.in_0_ready          (eth_tse_receive_ready),                     //         .ready
		.in_0_startofpacket  (eth_tse_receive_startofpacket),             //         .startofpacket
		.in_0_endofpacket    (eth_tse_receive_endofpacket),               //         .endofpacket
		.in_0_empty          (eth_tse_receive_empty),                     //         .empty
		.in_0_error          (eth_tse_receive_error),                     //         .error
		.out_0_data          (avalon_st_adapter_001_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_001_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_001_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_001_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_001_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_001_out_0_empty),         //         .empty
		.out_0_error         (avalon_st_adapter_001_out_0_error)          //         .error
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~mem_resetn_in_reset_reset_n),   // reset_in0.reset
		.clk            (sys_clk_clk),                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (sys_clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (cpu_debug_reset_request_reset),      // reset_in0.reset
		.reset_in1      (~mem_resetn_in_reset_reset_n),       // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (cpu_debug_reset_request_reset),      // reset_in0.reset
		.reset_in1      (~mem_resetn_in_reset_reset_n),       // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),          // reset_in1.reset
		.clk            (sys_clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_004_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_005 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (clock_bridge_0_in_clk_clk),          //       clk.clk
		.reset_out      (rst_controller_005_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_006 (
		.reset_in0      (cpu_debug_reset_request_reset),      // reset_in0.reset
		.reset_in1      (~mem_resetn_in_reset_reset_n),       // reset_in1.reset
		.clk            (ddr3_ram_afi_clk_clk),               //       clk.clk
		.reset_out      (rst_controller_006_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
