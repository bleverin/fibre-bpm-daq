// cali_ram.v

// Generated using ACDS version 19.1 670

`timescale 1 ps / 1 ps
module cali_ram (
		input  wire        cali_ram_clk1_clk,      //   cali_ram_clk1.clk
		input  wire        cali_ram_clk2_clk,      //   cali_ram_clk2.clk
		input  wire        cali_ram_reset1_reset,  // cali_ram_reset1.reset
		input  wire        cali_ram_reset2_reset,  // cali_ram_reset2.reset
		input  wire [8:0]  cali_ram_s1_address,    //     cali_ram_s1.address
		input  wire        cali_ram_s1_clken,      //                .clken
		input  wire        cali_ram_s1_chipselect, //                .chipselect
		input  wire        cali_ram_s1_write,      //                .write
		output wire [15:0] cali_ram_s1_readdata,   //                .readdata
		input  wire [15:0] cali_ram_s1_writedata,  //                .writedata
		input  wire [1:0]  cali_ram_s1_byteenable, //                .byteenable
		input  wire [8:0]  cali_ram_s2_address,    //     cali_ram_s2.address
		input  wire        cali_ram_s2_chipselect, //                .chipselect
		input  wire        cali_ram_s2_clken,      //                .clken
		input  wire        cali_ram_s2_write,      //                .write
		output wire [15:0] cali_ram_s2_readdata,   //                .readdata
		input  wire [15:0] cali_ram_s2_writedata,  //                .writedata
		input  wire [1:0]  cali_ram_s2_byteenable  //                .byteenable
	);

	cali_ram_cali_ram cali_ram (
		.clk         (cali_ram_clk1_clk),      //   clk1.clk
		.address     (cali_ram_s1_address),    //     s1.address
		.clken       (cali_ram_s1_clken),      //       .clken
		.chipselect  (cali_ram_s1_chipselect), //       .chipselect
		.write       (cali_ram_s1_write),      //       .write
		.readdata    (cali_ram_s1_readdata),   //       .readdata
		.writedata   (cali_ram_s1_writedata),  //       .writedata
		.byteenable  (cali_ram_s1_byteenable), //       .byteenable
		.reset       (cali_ram_reset1_reset),  // reset1.reset
		.address2    (cali_ram_s2_address),    //     s2.address
		.chipselect2 (cali_ram_s2_chipselect), //       .chipselect
		.clken2      (cali_ram_s2_clken),      //       .clken
		.write2      (cali_ram_s2_write),      //       .write
		.readdata2   (cali_ram_s2_readdata),   //       .readdata
		.writedata2  (cali_ram_s2_writedata),  //       .writedata
		.byteenable2 (cali_ram_s2_byteenable), //       .byteenable
		.clk2        (cali_ram_clk2_clk),      //   clk2.clk
		.reset2      (cali_ram_reset2_reset),  // reset2.reset
		.reset_req   (1'b0),                   // (terminated)
		.freeze      (1'b0),                   // (terminated)
		.reset_req2  (1'b0)                    // (terminated)
	);

endmodule
