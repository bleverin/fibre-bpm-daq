// q_sys_ext_flash_soft_asmiblock_instance_name.v

// Generated using ACDS version 19.1 670

`timescale 1 ps / 1 ps
module q_sys_ext_flash_soft_asmiblock_instance_name #(
		parameter IO_MODE  = "QUAD",
		parameter CS_WIDTH = 1
	) (
		input  wire       dclk,     //     dclk.conduit_dclk
		input  wire [0:0] sce,      //      sce.conduit_scein
		input  wire [3:0] dataout,  //  dataout.conduit_sdoin
		input  wire [3:0] dataoe,   //   dataoe.conduit_dataoe
		output wire [3:0] datain,   //   datain.conduit_dataout
		output wire       dclk_out, // dclk_out.conduit_dclk_out
		output wire [0:0] ncs       //      ncs.conduit_ncs
	);

	generate
		// If any of the display statements (or deliberately broken
		// instantiations) within this generate block triggers then this module
		// has been instantiated this module with a set of parameters different
		// from those it was generated for.  This will usually result in a
		// non-functioning system.
		if (IO_MODE != "QUAD")
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					io_mode_check ( .error(1'b1) );
		end
		if (CS_WIDTH != 1)
		begin
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
			instantiated_with_wrong_parameters_error_see_comment_above
					cs_width_check ( .error(1'b1) );
		end
	endgenerate

	soft_asmiblock #(
		.IO_MODE  ("QUAD"),
		.CS_WIDTH (1)
	) soft_asmiblock_instance_name (
		.dclk     (dclk),     //     dclk.conduit_dclk
		.sce      (sce),      //      sce.conduit_scein
		.dataout  (dataout),  //  dataout.conduit_sdoin
		.dataoe   (dataoe),   //   dataoe.conduit_dataoe
		.datain   (datain),   //   datain.conduit_dataout
		.dclk_out (dclk_out), // dclk_out.conduit_dclk_out
		.ncs      (ncs)       //      ncs.conduit_ncs
	);

endmodule
