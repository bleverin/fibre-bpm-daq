//bkg_subtraction_pipe_tb.v

//testbench for bkg_subtraction_pipe

`timescale 1 ns / 1 ns
module bkg_subtraction_pipe_tb();

	localparam CLK_PERIOD = 20; 

	reg clk;
	reg rst;
	
	//avalon ST(Streaming) sink: 0 readlatency and 0 readallowence
	reg [31:0] data_in_data;
	wire 		  data_in_ready;
	wire		  data_in_valid;
	reg [1:0]  data_in_empty;
	reg		  data_in_startofpacket;
	wire		  data_in_endofpacket;
	
	//avalon ST(Streaming) source: 0 readlatency and 0 readallowence
	wire [31:0] data_out_data;          // data_out.data
	wire        data_out_empty;         //         .empty
	wire        data_out_endofpacket;   //         .endofpacket
	wire        data_out_startofpacket; //         .startofpacket
	reg         data_out_ready;         //         .ready
	wire        data_out_valid;          //         .valid

	reg [1:0] state;
	localparam STATE_IDLE = 2'd0;
	localparam STATE_SEND = 2'd1;
	localparam STATE_LOC = 2'd3;
	
	reg [7:0]	tx_ctr; //counter for how many data has been sent
	localparam WORDS_TO_SEND = 163;
	
	bkg_subtraction_pipe #(.BKG_FRAME(4)) bkg_subtraction_dut(
	
		.clk		(clk),
		.rst		(rst),
		
		.data_in_data		(data_in_data),
		.data_in_ready		(data_in_ready),
		.data_in_valid		(data_in_valid),
		.data_in_empty		(data_in_empty),
		.data_in_startofpacket		(data_in_startofpacket),
		.data_in_endofpacket			(data_in_endofpacket),
		
		.data_out_data		(data_out_data),
		.data_out_empty	(data_out_empty),
		.data_out_endofpacket		(data_out_endofpacket),
		.data_out_startofpacket		(data_out_startofpacket),
		.data_out_ready	(data_out_ready),
		.data_out_valid	(data_out_valid),
		
		.to_udp_ready(1'b1)
		
	);
	
	initial begin
	
	clk = 1'b1;
	rst = 1'b1;
	
	//data_in_data = 32'hFFFFFFFF;
	data_in_data = 0;
	data_in_empty = 2'b0;
	data_in_startofpacket = 1'b0;
	//data_in_endofpacket = 1'b0;
	
	data_out_ready = 1'b0;
	
	state = STATE_IDLE;
	
	
	#(CLK_PERIOD*2);
	rst = 1'b0;
	
	//the next sink is ready..
	#(CLK_PERIOD*20);
	data_out_ready = 1'b1;
	
	#1; //make sure startofpacket and endofpacket start after clk rising edge
	
	repeat(8) begin
		/******one packet*******/
		//start packet
		#(CLK_PERIOD*2);
		data_in_startofpacket = 1'b1;
		//end packet
//		#(CLK_PERIOD*163*4);
//		data_in_endofpacket = 1'b1;
		#(CLK_PERIOD*500);
	end
	
	
	#(CLK_PERIOD*200); $stop;
	
	end
	
	
	//clk
	always #(CLK_PERIOD/2) clk = ~ clk;
	
	assign data_in_valid = (state == STATE_SEND || data_in_startofpacket || data_in_endofpacket)? 1'b1 : 1'b0;
	assign data_in_endofpacket = (state == STATE_SEND && tx_ctr == WORDS_TO_SEND -1)? 1'b1: 1'b0;
	always @(posedge clk) begin
		case(state)
		STATE_IDLE:
		begin
			tx_ctr <= 8'd0;
			if (data_in_startofpacket)
			begin
				state <= STATE_SEND;
				data_in_data <= data_in_data +1'b1;
			end
		end
		STATE_SEND:
		begin
			if (data_in_ready)
			begin
				data_in_startofpacket <= 1'b0;
				tx_ctr <= tx_ctr + 1'b1;
				if (tx_ctr == WORDS_TO_SEND-1) begin
					state <= STATE_LOC;
					data_in_data = 0;

					//data_in_data <= 32'hFFFFFFFF;
					//data_in_endofpacket <= 1'b0;
				end else begin
					data_in_data <= data_in_data +1'b1;
				end
			end
		end
		STATE_LOC:
		begin
			state <= STATE_IDLE;
			tx_ctr <= 8'd0;
		end
		endcase
	end
	
endmodule	