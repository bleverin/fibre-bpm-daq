
module sensor_algo (
	);	

endmodule
