// sensor_recon.v

// Generated using ACDS version 19.1 670

`timescale 1 ps / 1 ps
module sensor_recon (
		output wire [8:0]  sensor_recon_0_calibration_ram_interface_address,     // sensor_recon_0_calibration_ram_interface.address
		output wire        sensor_recon_0_calibration_ram_interface_read,        //                                         .read
		input  wire [15:0] sensor_recon_0_calibration_ram_interface_readdata,    //                                         .readdata
		input  wire        sensor_recon_0_calibration_ram_interface_waitrequest, //                                         .waitrequest
		input  wire        sensor_recon_0_clk_clk,                               //                       sensor_recon_0_clk.clk
		input  wire [1:0]  sensor_recon_0_csr_address,                           //                       sensor_recon_0_csr.address
		input  wire        sensor_recon_0_csr_read,                              //                                         .read
		output wire [31:0] sensor_recon_0_csr_readdata,                          //                                         .readdata
		input  wire        sensor_recon_0_csr_write,                             //                                         .write
		input  wire [31:0] sensor_recon_0_csr_writedata,                         //                                         .writedata
		input  wire [3:0]  sensor_recon_0_csr_byteenable,                        //                                         .byteenable
		output wire        sensor_recon_0_data_out_endofpacket,                  //                  sensor_recon_0_data_out.endofpacket
		output wire [31:0] sensor_recon_0_data_out_data,                         //                                         .data
		output wire [1:0]  sensor_recon_0_data_out_empty,                        //                                         .empty
		input  wire        sensor_recon_0_data_out_ready,                        //                                         .ready
		output wire        sensor_recon_0_data_out_startofpacket,                //                                         .startofpacket
		output wire        sensor_recon_0_data_out_valid,                        //                                         .valid
		input  wire        sensor_recon_0_rst_reset,                             //                       sensor_recon_0_rst.reset
		input  wire [4:0]  sensor_recon_0_sensor_in_adc_data,                    //                    sensor_recon_0_sensor.in_adc_data
		input  wire        sensor_recon_0_sensor_in_trg,                         //                                         .in_trg
		output wire        sensor_recon_0_sensor_out_adc_clk,                    //                                         .out_adc_clk
		output wire        sensor_recon_0_sensor_out_adc_cnv,                    //                                         .out_adc_cnv
		output wire        sensor_recon_0_sensor_out_sensor_clk,                 //                                         .out_sensor_clk
		output wire        sensor_recon_0_sensor_out_sensor_gain,                //                                         .out_sensor_gain
		output wire        sensor_recon_0_sensor_out_sensor_rst,                 //                                         .out_sensor_rst
		output wire [7:0]  sensor_recon_0_status_out_status_out,                 //                sensor_recon_0_status_out.status_out
		input  wire [7:0]  sensor_recon_0_synchro_ext_input,                     //                   sensor_recon_0_synchro.ext_input
		input  wire        sensor_recon_0_synchro_serial_rx,                     //                                         .serial_rx
		output wire        sensor_recon_0_synchro_serial_tx                      //                                         .serial_tx
	);

	sensor_algo sensor_recon_0 (
		.csr_address            (sensor_recon_0_csr_address),                           //                       csr.address
		.csr_read               (sensor_recon_0_csr_read),                              //                          .read
		.csr_readdata           (sensor_recon_0_csr_readdata),                          //                          .readdata
		.csr_write              (sensor_recon_0_csr_write),                             //                          .write
		.csr_writedata          (sensor_recon_0_csr_writedata),                         //                          .writedata
		.csr_byteenable         (sensor_recon_0_csr_byteenable),                        //                          .byteenable
		.data_out_endofpacket   (sensor_recon_0_data_out_endofpacket),                  //                  data_out.endofpacket
		.data_out_data          (sensor_recon_0_data_out_data),                         //                          .data
		.data_out_empty         (sensor_recon_0_data_out_empty),                        //                          .empty
		.data_out_ready         (sensor_recon_0_data_out_ready),                        //                          .ready
		.data_out_startofpacket (sensor_recon_0_data_out_startofpacket),                //                          .startofpacket
		.data_out_valid         (sensor_recon_0_data_out_valid),                        //                          .valid
		.clk_clk                (sensor_recon_0_clk_clk),                               //                       clk.clk
		.rst_reset              (sensor_recon_0_rst_reset),                             //                       rst.reset
		.in_adc_data            (sensor_recon_0_sensor_in_adc_data),                    //                    sensor.in_adc_data
		.in_trg                 (sensor_recon_0_sensor_in_trg),                         //                          .in_trg
		.out_adc_clk            (sensor_recon_0_sensor_out_adc_clk),                    //                          .out_adc_clk
		.out_adc_cnv            (sensor_recon_0_sensor_out_adc_cnv),                    //                          .out_adc_cnv
		.out_sensor_clk         (sensor_recon_0_sensor_out_sensor_clk),                 //                          .out_sensor_clk
		.out_sensor_gain        (sensor_recon_0_sensor_out_sensor_gain),                //                          .out_sensor_gain
		.out_sensor_rst         (sensor_recon_0_sensor_out_sensor_rst),                 //                          .out_sensor_rst
		.status_out             (sensor_recon_0_status_out_status_out),                 //                status_out.status_out
		.ext_input              (sensor_recon_0_synchro_ext_input),                     //                   synchro.ext_input
		.serial_rx              (sensor_recon_0_synchro_serial_rx),                     //                          .serial_rx
		.serial_tx              (sensor_recon_0_synchro_serial_tx),                     //                          .serial_tx
		.address                (sensor_recon_0_calibration_ram_interface_address),     // calibration_ram_interface.address
		.clken                  (sensor_recon_0_calibration_ram_interface_read),        //                          .read
		.cali_fac               (sensor_recon_0_calibration_ram_interface_readdata),    //                          .readdata
		.waitrequest            (sensor_recon_0_calibration_ram_interface_waitrequest)  //                          .waitrequest
	);

endmodule
