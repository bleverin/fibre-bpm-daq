// sensor_algo.v

// Generated using ACDS version 19.1 670

`timescale 1 ps / 1 ps
module sensor_algo (
		input  wire  sensor_algo_0_clk_clk,   // sensor_algo_0_clk.clk
		input  wire  sensor_algo_0_rst_reset  // sensor_algo_0_rst.reset
	);

	sensor_algo sensor_algo_0 (
		.csr_address            (),                        //           csr.address
		.csr_read               (),                        //              .read
		.csr_readdata           (),                        //              .readdata
		.csr_write              (),                        //              .write
		.csr_writedata          (),                        //              .writedata
		.csr_byteenable         (),                        //              .byteenable
		.clk_clk                (sensor_algo_0_clk_clk),   //           clk.clk
		.rst_reset              (sensor_algo_0_rst_reset), //           rst.reset
		.data_out_data          (),                        //      data_out.data
		.data_out_empty         (),                        //              .empty
		.data_out_ready         (),                        //              .ready
		.data_out_startofpacket (),                        //              .startofpacket
		.data_out_valid         (),                        //              .valid
		.data_out_endofpacket   (),                        //              .endofpacket
		.in_adc_data            (),                        //        sensor.in_adc_data
		.in_trg                 (),                        //              .in_trg
		.out_adc_clk            (),                        //              .out_adc_clk
		.out_adc_cnv            (),                        //              .out_adc_cnv
		.out_sensor_clk         (),                        //              .out_sensor_clk
		.out_sensor_gain        (),                        //              .out_sensor_gain
		.out_sensor_rst         (),                        //              .out_sensor_rst
		.ext_input              (),                        //       synchro.ext_input
		.serial_rx              (),                        //              .serial_rx
		.serial_tx              (),                        //              .serial_tx
		.status_out             (),                        //    status_out.status_out
		.address                (),                        // avalon_master.address
		.clken                  (),                        //              .read
		.cali_fac               ()                         //              .readdata
	);

endmodule
